// This is the unpowered netlist.
module divider (clk,
    cout1,
    cout10,
    cout2,
    cout3,
    cout4,
    cout5,
    cout6,
    cout7,
    cout8,
    cout9);
 input clk;
 output cout1;
 output cout10;
 output cout2;
 output cout3;
 output cout4;
 output cout5;
 output cout6;
 output cout7;
 output cout8;
 output cout9;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire clknet_leaf_0_clk;
 wire net235;
 wire net234;
 wire net233;
 wire net232;
 wire net231;
 wire net230;
 wire net229;
 wire net228;
 wire net227;
 wire net226;
 wire net225;
 wire net224;
 wire net223;
 wire net222;
 wire net221;
 wire net220;
 wire net219;
 wire net218;
 wire net217;
 wire net216;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire net215;
 wire net214;
 wire net213;
 wire net212;
 wire net211;
 wire net210;
 wire net209;
 wire net208;
 wire net207;
 wire net206;
 wire net205;
 wire net204;
 wire net203;
 wire net202;
 wire net201;
 wire net200;
 wire net199;
 wire net198;
 wire net197;
 wire net196;
 wire net195;
 wire net194;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire net193;
 wire net192;
 wire net191;
 wire net190;
 wire net189;
 wire net188;
 wire net187;
 wire net186;
 wire net185;
 wire net184;
 wire net183;
 wire net182;
 wire net181;
 wire net180;
 wire net179;
 wire net178;
 wire net177;
 wire net176;
 wire net175;
 wire net174;
 wire net173;
 wire net172;
 wire net171;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire net170;
 wire net169;
 wire net168;
 wire net167;
 wire net166;
 wire net165;
 wire net164;
 wire net163;
 wire net162;
 wire net161;
 wire net160;
 wire net159;
 wire net158;
 wire net157;
 wire net156;
 wire net155;
 wire net154;
 wire net153;
 wire net152;
 wire net151;
 wire net150;
 wire net149;
 wire net148;
 wire net147;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire net146;
 wire net145;
 wire net144;
 wire net143;
 wire net142;
 wire net141;
 wire net140;
 wire net139;
 wire net138;
 wire net137;
 wire net136;
 wire net135;
 wire net134;
 wire net133;
 wire net132;
 wire net131;
 wire net130;
 wire net129;
 wire net128;
 wire net127;
 wire net126;
 wire net125;
 wire net124;
 wire net123;
 wire net122;
 wire _0149_;
 wire _0150_;
 wire net121;
 wire net120;
 wire net119;
 wire net118;
 wire net117;
 wire net116;
 wire net115;
 wire net114;
 wire net113;
 wire net112;
 wire net111;
 wire net110;
 wire net109;
 wire net108;
 wire net107;
 wire net106;
 wire net105;
 wire net104;
 wire net103;
 wire net102;
 wire net101;
 wire net100;
 wire net99;
 wire net98;
 wire net97;
 wire net96;
 wire _0177_;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire net68;
 wire net67;
 wire net66;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire \counter10[0] ;
 wire \counter10[10] ;
 wire \counter10[11] ;
 wire \counter10[12] ;
 wire \counter10[13] ;
 wire \counter10[14] ;
 wire \counter10[15] ;
 wire \counter10[16] ;
 wire \counter10[17] ;
 wire \counter10[18] ;
 wire \counter10[19] ;
 wire \counter10[1] ;
 wire \counter10[20] ;
 wire \counter10[21] ;
 wire \counter10[22] ;
 wire \counter10[23] ;
 wire \counter10[24] ;
 wire \counter10[25] ;
 wire \counter10[26] ;
 wire \counter10[27] ;
 wire \counter10[2] ;
 wire \counter10[3] ;
 wire \counter10[4] ;
 wire \counter10[5] ;
 wire \counter10[6] ;
 wire \counter10[7] ;
 wire \counter10[8] ;
 wire \counter10[9] ;
 wire \counter2[0] ;
 wire \counter2[10] ;
 wire \counter2[11] ;
 wire \counter2[12] ;
 wire \counter2[13] ;
 wire \counter2[14] ;
 wire \counter2[15] ;
 wire \counter2[16] ;
 wire \counter2[17] ;
 wire \counter2[18] ;
 wire \counter2[19] ;
 wire \counter2[1] ;
 wire \counter2[20] ;
 wire \counter2[21] ;
 wire \counter2[22] ;
 wire \counter2[23] ;
 wire \counter2[24] ;
 wire \counter2[25] ;
 wire \counter2[26] ;
 wire \counter2[27] ;
 wire \counter2[2] ;
 wire \counter2[3] ;
 wire \counter2[4] ;
 wire \counter2[5] ;
 wire \counter2[6] ;
 wire \counter2[7] ;
 wire \counter2[8] ;
 wire \counter2[9] ;
 wire \counter3[0] ;
 wire \counter3[10] ;
 wire \counter3[11] ;
 wire \counter3[12] ;
 wire \counter3[13] ;
 wire \counter3[14] ;
 wire \counter3[15] ;
 wire \counter3[16] ;
 wire \counter3[17] ;
 wire \counter3[18] ;
 wire \counter3[19] ;
 wire \counter3[1] ;
 wire \counter3[20] ;
 wire \counter3[21] ;
 wire \counter3[22] ;
 wire \counter3[23] ;
 wire \counter3[24] ;
 wire \counter3[25] ;
 wire \counter3[26] ;
 wire \counter3[27] ;
 wire \counter3[2] ;
 wire \counter3[3] ;
 wire \counter3[4] ;
 wire \counter3[5] ;
 wire \counter3[6] ;
 wire \counter3[7] ;
 wire \counter3[8] ;
 wire \counter3[9] ;
 wire \counter4[0] ;
 wire \counter4[10] ;
 wire \counter4[11] ;
 wire \counter4[12] ;
 wire \counter4[13] ;
 wire \counter4[14] ;
 wire \counter4[15] ;
 wire \counter4[16] ;
 wire \counter4[17] ;
 wire \counter4[18] ;
 wire \counter4[19] ;
 wire \counter4[1] ;
 wire \counter4[20] ;
 wire \counter4[21] ;
 wire \counter4[22] ;
 wire \counter4[23] ;
 wire \counter4[24] ;
 wire \counter4[25] ;
 wire \counter4[26] ;
 wire \counter4[27] ;
 wire \counter4[2] ;
 wire \counter4[3] ;
 wire \counter4[4] ;
 wire \counter4[5] ;
 wire \counter4[6] ;
 wire \counter4[7] ;
 wire \counter4[8] ;
 wire \counter4[9] ;
 wire \counter5[0] ;
 wire \counter5[10] ;
 wire \counter5[11] ;
 wire \counter5[12] ;
 wire \counter5[13] ;
 wire \counter5[14] ;
 wire \counter5[15] ;
 wire \counter5[16] ;
 wire \counter5[17] ;
 wire \counter5[18] ;
 wire \counter5[19] ;
 wire \counter5[1] ;
 wire \counter5[20] ;
 wire \counter5[21] ;
 wire \counter5[22] ;
 wire \counter5[23] ;
 wire \counter5[24] ;
 wire \counter5[25] ;
 wire \counter5[26] ;
 wire \counter5[27] ;
 wire \counter5[2] ;
 wire \counter5[3] ;
 wire \counter5[4] ;
 wire \counter5[5] ;
 wire \counter5[6] ;
 wire \counter5[7] ;
 wire \counter5[8] ;
 wire \counter5[9] ;
 wire \counter6[0] ;
 wire \counter6[10] ;
 wire \counter6[11] ;
 wire \counter6[12] ;
 wire \counter6[13] ;
 wire \counter6[14] ;
 wire \counter6[15] ;
 wire \counter6[16] ;
 wire \counter6[17] ;
 wire \counter6[18] ;
 wire \counter6[19] ;
 wire \counter6[1] ;
 wire \counter6[20] ;
 wire \counter6[21] ;
 wire \counter6[22] ;
 wire \counter6[23] ;
 wire \counter6[24] ;
 wire \counter6[25] ;
 wire \counter6[26] ;
 wire \counter6[27] ;
 wire \counter6[2] ;
 wire \counter6[3] ;
 wire \counter6[4] ;
 wire \counter6[5] ;
 wire \counter6[6] ;
 wire \counter6[7] ;
 wire \counter6[8] ;
 wire \counter6[9] ;
 wire \counter7[0] ;
 wire \counter7[10] ;
 wire \counter7[11] ;
 wire \counter7[12] ;
 wire \counter7[13] ;
 wire \counter7[14] ;
 wire \counter7[15] ;
 wire \counter7[16] ;
 wire \counter7[17] ;
 wire \counter7[18] ;
 wire \counter7[19] ;
 wire \counter7[1] ;
 wire \counter7[20] ;
 wire \counter7[21] ;
 wire \counter7[22] ;
 wire \counter7[23] ;
 wire \counter7[24] ;
 wire \counter7[25] ;
 wire \counter7[26] ;
 wire \counter7[27] ;
 wire \counter7[2] ;
 wire \counter7[3] ;
 wire \counter7[4] ;
 wire \counter7[5] ;
 wire \counter7[6] ;
 wire \counter7[7] ;
 wire \counter7[8] ;
 wire \counter7[9] ;
 wire \counter8[0] ;
 wire \counter8[10] ;
 wire \counter8[11] ;
 wire \counter8[12] ;
 wire \counter8[13] ;
 wire \counter8[14] ;
 wire \counter8[15] ;
 wire \counter8[16] ;
 wire \counter8[17] ;
 wire \counter8[18] ;
 wire \counter8[19] ;
 wire \counter8[1] ;
 wire \counter8[20] ;
 wire \counter8[21] ;
 wire \counter8[22] ;
 wire \counter8[23] ;
 wire \counter8[24] ;
 wire \counter8[25] ;
 wire \counter8[26] ;
 wire \counter8[27] ;
 wire \counter8[2] ;
 wire \counter8[3] ;
 wire \counter8[4] ;
 wire \counter8[5] ;
 wire \counter8[6] ;
 wire \counter8[7] ;
 wire \counter8[8] ;
 wire \counter8[9] ;
 wire \counter9[0] ;
 wire \counter9[10] ;
 wire \counter9[11] ;
 wire \counter9[12] ;
 wire \counter9[13] ;
 wire \counter9[14] ;
 wire \counter9[15] ;
 wire \counter9[16] ;
 wire \counter9[17] ;
 wire \counter9[18] ;
 wire \counter9[19] ;
 wire \counter9[1] ;
 wire \counter9[20] ;
 wire \counter9[21] ;
 wire \counter9[22] ;
 wire \counter9[23] ;
 wire \counter9[24] ;
 wire \counter9[25] ;
 wire \counter9[26] ;
 wire \counter9[27] ;
 wire \counter9[2] ;
 wire \counter9[3] ;
 wire \counter9[4] ;
 wire \counter9[5] ;
 wire \counter9[6] ;
 wire \counter9[7] ;
 wire \counter9[8] ;
 wire \counter9[9] ;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[16] ;
 wire \counter[17] ;
 wire \counter[18] ;
 wire \counter[19] ;
 wire \counter[1] ;
 wire \counter[20] ;
 wire \counter[21] ;
 wire \counter[22] ;
 wire \counter[23] ;
 wire \counter[24] ;
 wire \counter[25] ;
 wire \counter[26] ;
 wire \counter[27] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0475_ (.A1(\counter[20] ),
    .A2(\counter[19] ),
    .A3(\counter[18] ),
    .A4(\counter[17] ),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0476_ (.A1(\counter[16] ),
    .A2(\counter[15] ),
    .A3(\counter[13] ),
    .A4(\counter[14] ),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0477_ (.A1(\counter[24] ),
    .A2(\counter[23] ),
    .A3(\counter[22] ),
    .A4(\counter[21] ),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0478_ (.A1(\counter[26] ),
    .A2(\counter[25] ),
    .A3(\counter[1] ),
    .A4(\counter[0] ),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0479_ (.A1(_0306_),
    .A2(_0307_),
    .A3(_0308_),
    .A4(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0480_ (.A1(\counter[4] ),
    .A2(\counter[3] ),
    .A3(\counter[2] ),
    .A4(\counter[27] ),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0481_ (.A1(\counter[8] ),
    .A2(\counter[7] ),
    .A3(\counter[6] ),
    .A4(\counter[5] ),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0482_ (.A1(\counter[12] ),
    .A2(\counter[11] ),
    .A3(\counter[9] ),
    .A4(\counter[10] ),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0483_ (.A1(_0311_),
    .A2(_0312_),
    .A3(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0484_ (.A1(_0310_),
    .A2(_0314_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0485_ (.A1(\counter2[5] ),
    .A2(\counter2[4] ),
    .A3(\counter2[3] ),
    .A4(\counter2[2] ),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0486_ (.A1(\counter2[9] ),
    .A2(\counter2[8] ),
    .A3(\counter2[7] ),
    .A4(\counter2[6] ),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0487_ (.A1(\counter2[13] ),
    .A2(\counter2[12] ),
    .A3(\counter2[11] ),
    .A4(\counter2[10] ),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0488_ (.A1(\counter2[1] ),
    .A2(\counter2[0] ),
    .B(\counter2[27] ),
    .C(\counter2[26] ),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0489_ (.A1(\counter2[25] ),
    .A2(\counter2[24] ),
    .A3(\counter2[23] ),
    .A4(\counter2[22] ),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0490_ (.A1(\counter2[21] ),
    .A2(\counter2[20] ),
    .A3(\counter2[19] ),
    .A4(\counter2[18] ),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0491_ (.A1(\counter2[17] ),
    .A2(\counter2[16] ),
    .A3(\counter2[15] ),
    .A4(\counter2[14] ),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0492_ (.A1(_0318_),
    .A2(_0319_),
    .A3(_0320_),
    .A4(_0321_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0493_ (.A1(_0315_),
    .A2(_0316_),
    .A3(_0317_),
    .A4(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0494_ (.A1(\counter2[1] ),
    .A2(_0323_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0495_ (.A1(\counter3[4] ),
    .A2(\counter3[3] ),
    .A3(\counter3[27] ),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0496_ (.A1(\counter3[7] ),
    .A2(\counter3[8] ),
    .A3(\counter3[6] ),
    .A4(\counter3[5] ),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0497_ (.A1(\counter3[12] ),
    .A2(\counter3[11] ),
    .A3(\counter3[10] ),
    .A4(\counter3[9] ),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0498_ (.A1(\counter3[25] ),
    .A2(\counter3[26] ),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0499_ (.A1(\counter3[24] ),
    .A2(\counter3[23] ),
    .A3(\counter3[22] ),
    .A4(\counter3[21] ),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0500_ (.A1(\counter3[20] ),
    .A2(\counter3[19] ),
    .A3(\counter3[18] ),
    .A4(\counter3[17] ),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0501_ (.A1(\counter3[16] ),
    .A2(\counter3[15] ),
    .A3(\counter3[14] ),
    .A4(\counter3[13] ),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0502_ (.A1(_0327_),
    .A2(_0328_),
    .A3(_0329_),
    .A4(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0503_ (.A1(_0324_),
    .A2(_0325_),
    .A3(_0326_),
    .A4(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0504_ (.A1(\counter3[2] ),
    .A2(_0332_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0505_ (.A1(\counter4[22] ),
    .A2(\counter4[23] ),
    .A3(\counter4[21] ),
    .A4(\counter4[20] ),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0506_ (.A1(\counter4[27] ),
    .A2(\counter4[26] ),
    .A3(\counter4[24] ),
    .A4(\counter4[25] ),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0507_ (.A1(\counter4[14] ),
    .A2(\counter4[15] ),
    .A3(\counter4[12] ),
    .A4(\counter4[13] ),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0508_ (.A1(\counter4[18] ),
    .A2(\counter4[19] ),
    .A3(\counter4[17] ),
    .A4(\counter4[16] ),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0509_ (.A1(\counter4[11] ),
    .A2(\counter4[10] ),
    .A3(\counter4[9] ),
    .A4(\counter4[8] ),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0510_ (.A1(\counter4[7] ),
    .A2(\counter4[6] ),
    .A3(\counter4[5] ),
    .A4(\counter4[4] ),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0511_ (.A1(_0335_),
    .A2(_0336_),
    .A3(_0337_),
    .A4(_0338_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0512_ (.A1(_0333_),
    .A2(_0334_),
    .A3(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0513_ (.I(_0340_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0514_ (.A1(\counter4[3] ),
    .A2(_0341_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0515_ (.A1(\counter5[22] ),
    .A2(\counter5[21] ),
    .A3(\counter5[20] ),
    .A4(\counter5[19] ),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0516_ (.A1(\counter5[26] ),
    .A2(\counter5[25] ),
    .A3(\counter5[24] ),
    .A4(\counter5[23] ),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0517_ (.A1(\counter5[14] ),
    .A2(\counter5[13] ),
    .A3(\counter5[12] ),
    .A4(\counter5[11] ),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0518_ (.A1(\counter5[18] ),
    .A2(\counter5[17] ),
    .A3(\counter5[16] ),
    .A4(\counter5[15] ),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0519_ (.A1(\counter5[10] ),
    .A2(\counter5[9] ),
    .A3(\counter5[8] ),
    .A4(\counter5[7] ),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0520_ (.A1(\counter5[6] ),
    .A2(\counter5[5] ),
    .A3(\counter5[27] ),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0521_ (.A1(_0344_),
    .A2(_0345_),
    .A3(_0346_),
    .A4(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0522_ (.A1(_0342_),
    .A2(_0343_),
    .A3(_0348_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0523_ (.I(_0349_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0524_ (.A1(\counter5[4] ),
    .A2(_0350_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0525_ (.A1(\counter6[25] ),
    .A2(\counter6[24] ),
    .A3(\counter6[23] ),
    .A4(\counter6[22] ),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0526_ (.A1(\counter6[27] ),
    .A2(\counter6[26] ),
    .A3(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0527_ (.A1(\counter6[17] ),
    .A2(\counter6[16] ),
    .A3(\counter6[14] ),
    .A4(\counter6[15] ),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0528_ (.A1(\counter6[21] ),
    .A2(\counter6[20] ),
    .A3(\counter6[18] ),
    .A4(\counter6[19] ),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0529_ (.A1(_0353_),
    .A2(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0530_ (.A1(\counter6[13] ),
    .A2(\counter6[12] ),
    .A3(\counter6[10] ),
    .A4(\counter6[11] ),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0531_ (.A1(\counter6[9] ),
    .A2(\counter6[8] ),
    .A3(\counter6[7] ),
    .A4(\counter6[6] ),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0532_ (.A1(_0356_),
    .A2(_0357_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0533_ (.A1(_0352_),
    .A2(_0355_),
    .A3(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0534_ (.A1(\counter6[5] ),
    .A2(_0359_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0535_ (.A1(\counter7[27] ),
    .A2(\counter7[26] ),
    .A3(\counter7[7] ),
    .A4(\counter7[8] ),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0536_ (.A1(\counter7[25] ),
    .A2(\counter7[24] ),
    .A3(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0537_ (.A1(\counter7[13] ),
    .A2(\counter7[14] ),
    .A3(\counter7[15] ),
    .A4(\counter7[16] ),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0538_ (.A1(\counter7[9] ),
    .A2(\counter7[10] ),
    .A3(\counter7[11] ),
    .A4(\counter7[12] ),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0539_ (.A1(_0362_),
    .A2(_0363_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0540_ (.A1(\counter7[17] ),
    .A2(\counter7[18] ),
    .A3(\counter7[19] ),
    .A4(\counter7[20] ),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0541_ (.A1(\counter7[21] ),
    .A2(\counter7[22] ),
    .A3(\counter7[23] ),
    .A4(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0542_ (.A1(_0361_),
    .A2(_0364_),
    .A3(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0543_ (.A1(\counter7[6] ),
    .A2(_0367_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0544_ (.A1(\counter8[20] ),
    .A2(\counter8[21] ),
    .A3(\counter8[23] ),
    .A4(\counter8[22] ),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0545_ (.A1(\counter8[27] ),
    .A2(\counter8[26] ),
    .A3(\counter8[24] ),
    .A4(\counter8[25] ),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0546_ (.A1(_0368_),
    .A2(_0369_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0547_ (.A1(\counter8[10] ),
    .A2(\counter8[11] ),
    .A3(\counter8[9] ),
    .A4(\counter8[8] ),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0548_ (.A1(\counter8[12] ),
    .A2(\counter8[13] ),
    .A3(\counter8[14] ),
    .A4(\counter8[15] ),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0549_ (.A1(\counter8[18] ),
    .A2(\counter8[19] ),
    .A3(\counter8[17] ),
    .A4(\counter8[16] ),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0550_ (.A1(_0371_),
    .A2(_0372_),
    .A3(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0551_ (.A1(_0370_),
    .A2(_0374_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0552_ (.A1(\counter8[7] ),
    .A2(_0375_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0553_ (.I(\counter9[8] ),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0554_ (.A1(\counter9[22] ),
    .A2(\counter9[21] ),
    .A3(\counter9[20] ),
    .A4(\counter9[19] ),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0555_ (.A1(\counter9[26] ),
    .A2(\counter9[25] ),
    .A3(\counter9[23] ),
    .A4(\counter9[24] ),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0556_ (.A1(_0377_),
    .A2(_0378_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0557_ (.A1(\counter9[10] ),
    .A2(\counter9[9] ),
    .A3(\counter9[27] ),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0558_ (.A1(\counter9[14] ),
    .A2(\counter9[13] ),
    .A3(\counter9[12] ),
    .A4(\counter9[11] ),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0559_ (.A1(\counter9[18] ),
    .A2(\counter9[17] ),
    .A3(\counter9[16] ),
    .A4(\counter9[15] ),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0560_ (.A1(_0380_),
    .A2(_0381_),
    .A3(_0382_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0561_ (.A1(_0376_),
    .A2(_0379_),
    .A3(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0562_ (.I(_0384_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0563_ (.I(\counter10[9] ),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0564_ (.A1(\counter10[25] ),
    .A2(\counter10[24] ),
    .A3(\counter10[23] ),
    .A4(\counter10[22] ),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0565_ (.A1(\counter10[27] ),
    .A2(\counter10[26] ),
    .A3(_0386_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0566_ (.A1(\counter10[13] ),
    .A2(\counter10[12] ),
    .A3(\counter10[11] ),
    .A4(\counter10[10] ),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0567_ (.A1(\counter10[17] ),
    .A2(\counter10[16] ),
    .A3(\counter10[15] ),
    .A4(\counter10[14] ),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0568_ (.A1(\counter10[21] ),
    .A2(\counter10[20] ),
    .A3(\counter10[19] ),
    .A4(\counter10[18] ),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0569_ (.A1(_0388_),
    .A2(_0389_),
    .A3(_0390_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0570_ (.A1(_0385_),
    .A2(_0387_),
    .A3(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0571_ (.I(_0392_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0572_ (.I(_0393_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0573_ (.A1(\counter7[0] ),
    .A2(\counter7[1] ),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0574_ (.A1(\counter7[0] ),
    .A2(\counter7[3] ),
    .A3(\counter7[2] ),
    .A4(\counter7[1] ),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0575_ (.A1(\counter7[6] ),
    .A2(\counter7[5] ),
    .A3(\counter7[4] ),
    .A4(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0576_ (.A1(_0361_),
    .A2(_0364_),
    .A3(_0366_),
    .A4(_0396_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0577_ (.I(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0578_ (.A1(\counter7[0] ),
    .A2(\counter7[1] ),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0579_ (.A1(_0394_),
    .A2(_0398_),
    .A3(_0399_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0580_ (.A1(\counter7[2] ),
    .A2(_0394_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0581_ (.A1(_0398_),
    .A2(_0400_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0582_ (.A1(\counter7[2] ),
    .A2(_0394_),
    .B(\counter7[3] ),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0583_ (.A1(_0395_),
    .A2(_0397_),
    .A3(_0401_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0584_ (.A1(\counter7[4] ),
    .A2(_0395_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0585_ (.A1(\counter7[4] ),
    .A2(_0395_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0586_ (.A1(_0367_),
    .A2(_0402_),
    .A3(_0403_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0587_ (.A1(\counter7[5] ),
    .A2(_0402_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0588_ (.A1(\counter7[5] ),
    .A2(_0402_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0589_ (.A1(_0367_),
    .A2(_0404_),
    .A3(_0405_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0590_ (.A1(\counter7[5] ),
    .A2(_0402_),
    .B(\counter7[6] ),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0591_ (.A1(_0398_),
    .A2(_0406_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0592_ (.A1(\counter6[1] ),
    .A2(\counter6[0] ),
    .A3(\counter6[2] ),
    .A4(\counter6[3] ),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0593_ (.A1(\counter6[5] ),
    .A2(\counter6[4] ),
    .A3(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0594_ (.A1(_0352_),
    .A2(_0355_),
    .A3(_0358_),
    .A4(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0595_ (.A1(\counter6[0] ),
    .A2(_0409_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0596_ (.A1(\counter6[1] ),
    .A2(\counter6[0] ),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0597_ (.A1(\counter6[1] ),
    .A2(\counter6[0] ),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0598_ (.A1(_0410_),
    .A2(_0409_),
    .A3(_0411_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0599_ (.A1(\counter6[2] ),
    .A2(_0410_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0600_ (.A1(_0409_),
    .A2(_0412_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0601_ (.A1(\counter6[2] ),
    .A2(_0410_),
    .B(\counter6[3] ),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0602_ (.A1(_0359_),
    .A2(_0407_),
    .A3(_0413_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0603_ (.A1(\counter6[4] ),
    .A2(_0407_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0604_ (.A1(\counter6[4] ),
    .A2(_0407_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0605_ (.A1(_0359_),
    .A2(_0414_),
    .A3(_0415_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0606_ (.A1(\counter6[5] ),
    .A2(_0414_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0607_ (.A1(_0409_),
    .A2(_0416_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0608_ (.A1(\counter5[1] ),
    .A2(\counter5[0] ),
    .A3(\counter5[2] ),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0609_ (.A1(\counter5[3] ),
    .A2(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0610_ (.A1(\counter5[4] ),
    .A2(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0611_ (.A1(\counter5[0] ),
    .A2(_0350_),
    .A3(_0419_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0612_ (.A1(\counter5[1] ),
    .A2(\counter5[0] ),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0613_ (.A1(\counter5[1] ),
    .A2(\counter5[0] ),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0614_ (.A1(_0350_),
    .A2(_0420_),
    .A3(_0421_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0615_ (.A1(\counter5[2] ),
    .A2(_0420_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0616_ (.A1(_0350_),
    .A2(_0417_),
    .A3(_0422_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0617_ (.A1(\counter5[3] ),
    .A2(_0417_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0618_ (.A1(_0349_),
    .A2(_0418_),
    .A3(_0423_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0619_ (.A1(\counter5[4] ),
    .A2(_0418_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0620_ (.A1(_0349_),
    .A2(_0419_),
    .A3(_0424_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0621_ (.A1(\counter4[0] ),
    .A2(_0341_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0622_ (.A1(\counter4[0] ),
    .A2(\counter4[1] ),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0623_ (.A1(\counter4[0] ),
    .A2(\counter4[1] ),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0624_ (.A1(_0341_),
    .A2(_0425_),
    .A3(_0426_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0625_ (.A1(\counter4[2] ),
    .A2(_0425_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0626_ (.A1(\counter4[2] ),
    .A2(_0425_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0627_ (.A1(_0341_),
    .A2(_0427_),
    .A3(_0428_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0628_ (.A1(\counter4[3] ),
    .A2(_0427_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0629_ (.A1(\counter4[3] ),
    .A2(_0427_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0630_ (.A1(_0340_),
    .A2(_0429_),
    .A3(_0430_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0631_ (.A1(\counter3[0] ),
    .A2(_0332_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0632_ (.A1(\counter3[1] ),
    .A2(\counter3[0] ),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0633_ (.A1(_0332_),
    .A2(_0431_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0634_ (.A1(\counter3[1] ),
    .A2(\counter3[0] ),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0635_ (.A1(\counter3[2] ),
    .A2(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0636_ (.A1(_0332_),
    .A2(_0433_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0637_ (.A1(\counter2[0] ),
    .A2(_0323_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0638_ (.A1(\counter2[1] ),
    .A2(\counter2[0] ),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0639_ (.A1(_0323_),
    .A2(_0434_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0640_ (.A1(_0310_),
    .A2(_0314_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0641_ (.I(\counter10[8] ),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0642_ (.A1(\counter10[1] ),
    .A2(\counter10[0] ),
    .A3(\counter10[3] ),
    .A4(\counter10[2] ),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0643_ (.A1(\counter10[5] ),
    .A2(\counter10[4] ),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0644_ (.A1(\counter10[7] ),
    .A2(\counter10[6] ),
    .A3(_0436_),
    .A4(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0645_ (.A1(_0435_),
    .A2(_0438_),
    .B(_0391_),
    .C(_0387_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0646_ (.I(_0439_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0647_ (.I(\counter10[0] ),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0648_ (.A1(_0393_),
    .A2(_0440_),
    .B(_0441_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0649_ (.A1(\counter10[1] ),
    .A2(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0650_ (.A1(_0393_),
    .A2(_0440_),
    .B(_0442_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0651_ (.I(_0439_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0652_ (.A1(\counter10[1] ),
    .A2(_0441_),
    .B(\counter10[2] ),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0653_ (.A1(\counter10[1] ),
    .A2(_0441_),
    .A3(\counter10[2] ),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0654_ (.A1(_0392_),
    .A2(_0443_),
    .B(_0444_),
    .C(_0445_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0655_ (.A1(\counter10[3] ),
    .A2(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0656_ (.I(_0436_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0657_ (.A1(_0392_),
    .A2(_0439_),
    .B(_0446_),
    .C(_0447_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0658_ (.I(_0392_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0659_ (.A1(\counter10[4] ),
    .A2(_0447_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0660_ (.A1(_0448_),
    .A2(_0440_),
    .B(_0449_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0661_ (.A1(\counter10[4] ),
    .A2(_0447_),
    .B(\counter10[5] ),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0662_ (.A1(_0447_),
    .A2(_0437_),
    .B1(_0439_),
    .B2(_0448_),
    .C(_0450_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0663_ (.A1(_0436_),
    .A2(_0437_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0664_ (.A1(\counter10[6] ),
    .A2(_0451_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0665_ (.A1(_0448_),
    .A2(_0440_),
    .B(_0452_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0666_ (.A1(\counter10[6] ),
    .A2(_0436_),
    .A3(_0437_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0667_ (.A1(\counter10[7] ),
    .A2(_0453_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0668_ (.A1(_0448_),
    .A2(_0443_),
    .B(_0454_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0669_ (.A1(_0435_),
    .A2(_0438_),
    .B(_0443_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0670_ (.A1(_0435_),
    .A2(_0438_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0671_ (.A1(_0385_),
    .A2(_0455_),
    .B1(_0443_),
    .B2(_0393_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0672_ (.I(\counter9[0] ),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0673_ (.A1(\counter9[3] ),
    .A2(\counter9[2] ),
    .A3(\counter9[1] ),
    .A4(\counter9[0] ),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0674_ (.A1(\counter9[5] ),
    .A2(\counter9[4] ),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0675_ (.A1(\counter9[7] ),
    .A2(\counter9[6] ),
    .A3(_0457_),
    .A4(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0676_ (.A1(_0376_),
    .A2(_0459_),
    .B(_0383_),
    .C(_0379_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0677_ (.I(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0678_ (.A1(_0456_),
    .A2(_0461_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0679_ (.A1(\counter9[1] ),
    .A2(_0456_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0680_ (.A1(_0461_),
    .A2(_0462_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0681_ (.A1(\counter9[2] ),
    .A2(\counter9[1] ),
    .A3(_0456_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0682_ (.I(_0460_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0683_ (.A1(\counter9[1] ),
    .A2(_0456_),
    .B(\counter9[2] ),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0684_ (.A1(_0463_),
    .A2(_0464_),
    .A3(_0465_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0685_ (.I(_0457_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0686_ (.A1(\counter9[3] ),
    .A2(_0463_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0687_ (.A1(_0466_),
    .A2(_0464_),
    .A3(_0467_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0688_ (.A1(\counter9[4] ),
    .A2(_0457_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0689_ (.A1(_0461_),
    .A2(_0468_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0690_ (.A1(\counter9[4] ),
    .A2(_0466_),
    .B(\counter9[5] ),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0691_ (.A1(_0466_),
    .A2(_0458_),
    .B(_0464_),
    .C(_0469_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0692_ (.A1(_0457_),
    .A2(_0458_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _0693_ (.A1(\counter9[6] ),
    .A2(_0470_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0694_ (.A1(_0464_),
    .A2(_0471_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0695_ (.I(\counter9[7] ),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0696_ (.A1(\counter9[6] ),
    .A2(_0466_),
    .A3(_0458_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0697_ (.A1(_0379_),
    .A2(_0383_),
    .A3(_0459_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0698_ (.A1(_0472_),
    .A2(_0473_),
    .B(_0474_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0699_ (.A1(_0376_),
    .A2(_0459_),
    .B(_0461_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0700_ (.I(\counter8[0] ),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0701_ (.I(\counter8[7] ),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0702_ (.A1(\counter8[2] ),
    .A2(\counter8[3] ),
    .A3(\counter8[1] ),
    .A4(\counter8[0] ),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0703_ (.A1(\counter8[6] ),
    .A2(\counter8[4] ),
    .A3(\counter8[5] ),
    .A4(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0704_ (.A1(_0291_),
    .A2(_0293_),
    .B(_0374_),
    .C(_0370_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0705_ (.I(_0294_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0706_ (.A1(_0290_),
    .A2(_0295_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0707_ (.A1(\counter8[1] ),
    .A2(_0290_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0708_ (.A1(_0295_),
    .A2(_0296_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0709_ (.A1(\counter8[2] ),
    .A2(\counter8[1] ),
    .A3(_0290_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0710_ (.A1(\counter8[1] ),
    .A2(_0290_),
    .B(\counter8[2] ),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0711_ (.A1(_0297_),
    .A2(_0294_),
    .A3(_0298_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0712_ (.I(_0292_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0713_ (.A1(\counter8[3] ),
    .A2(_0297_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0714_ (.A1(_0299_),
    .A2(_0294_),
    .A3(_0300_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _0715_ (.A1(\counter8[4] ),
    .A2(_0299_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0716_ (.A1(_0295_),
    .A2(_0301_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0717_ (.A1(\counter8[4] ),
    .A2(\counter8[5] ),
    .A3(_0299_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0718_ (.A1(\counter8[4] ),
    .A2(_0299_),
    .B(\counter8[5] ),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0719_ (.A1(_0302_),
    .A2(_0294_),
    .A3(_0303_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0720_ (.I(_0293_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0721_ (.A1(\counter8[6] ),
    .A2(_0302_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0722_ (.A1(_0375_),
    .A2(_0304_),
    .A3(_0305_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0723_ (.A1(_0291_),
    .A2(_0293_),
    .B(_0295_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0724_ (.A1(\counter7[0] ),
    .A2(_0398_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0725_ (.D(_0010_),
    .CLK(clknet_leaf_14_clk),
    .Q(\counter7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0726_ (.D(_0011_),
    .CLK(clknet_leaf_14_clk),
    .Q(\counter7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0727_ (.D(_0012_),
    .CLK(clknet_leaf_13_clk),
    .Q(\counter7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0728_ (.D(_0013_),
    .CLK(clknet_leaf_11_clk),
    .Q(\counter7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0729_ (.D(_0014_),
    .CLK(clknet_leaf_12_clk),
    .Q(\counter7[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0730_ (.D(_0015_),
    .CLK(clknet_leaf_12_clk),
    .Q(\counter7[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0731_ (.D(net235),
    .CLK(clknet_leaf_11_clk),
    .Q(\counter7[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0732_ (.D(net234),
    .CLK(clknet_leaf_11_clk),
    .Q(\counter7[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0733_ (.D(net233),
    .CLK(clknet_leaf_14_clk),
    .Q(\counter7[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0734_ (.D(net232),
    .CLK(clknet_leaf_13_clk),
    .Q(\counter7[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0735_ (.D(net231),
    .CLK(clknet_leaf_10_clk),
    .Q(\counter7[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0736_ (.D(net230),
    .CLK(clknet_leaf_10_clk),
    .Q(\counter7[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0737_ (.D(net229),
    .CLK(clknet_leaf_7_clk),
    .Q(\counter7[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0738_ (.D(net228),
    .CLK(clknet_leaf_7_clk),
    .Q(\counter7[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0739_ (.D(net227),
    .CLK(clknet_leaf_10_clk),
    .Q(\counter7[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0740_ (.D(net226),
    .CLK(clknet_leaf_9_clk),
    .Q(\counter7[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0741_ (.D(net225),
    .CLK(clknet_leaf_9_clk),
    .Q(\counter7[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0742_ (.D(net224),
    .CLK(clknet_leaf_9_clk),
    .Q(\counter7[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0743_ (.D(net223),
    .CLK(clknet_leaf_7_clk),
    .Q(\counter7[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0744_ (.D(net222),
    .CLK(clknet_leaf_8_clk),
    .Q(\counter7[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0745_ (.D(net221),
    .CLK(clknet_leaf_10_clk),
    .Q(\counter7[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0746_ (.D(net220),
    .CLK(clknet_leaf_9_clk),
    .Q(\counter7[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0747_ (.D(net219),
    .CLK(clknet_leaf_9_clk),
    .Q(\counter7[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0748_ (.D(net218),
    .CLK(clknet_leaf_10_clk),
    .Q(\counter7[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0749_ (.D(net217),
    .CLK(clknet_leaf_11_clk),
    .Q(\counter7[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0750_ (.D(net216),
    .CLK(clknet_leaf_11_clk),
    .Q(\counter7[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0751_ (.D(net215),
    .CLK(clknet_leaf_11_clk),
    .Q(\counter7[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0752_ (.D(_0005_),
    .CLK(clknet_leaf_25_clk),
    .Q(net6));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0753_ (.D(_0037_),
    .CLK(clknet_leaf_48_clk),
    .Q(\counter6[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0754_ (.D(_0038_),
    .CLK(clknet_leaf_41_clk),
    .Q(\counter6[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0755_ (.D(_0039_),
    .CLK(clknet_leaf_47_clk),
    .Q(\counter6[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0756_ (.D(_0040_),
    .CLK(clknet_leaf_48_clk),
    .Q(\counter6[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0757_ (.D(_0041_),
    .CLK(clknet_leaf_48_clk),
    .Q(\counter6[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0758_ (.D(_0042_),
    .CLK(clknet_leaf_48_clk),
    .Q(\counter6[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0759_ (.D(net214),
    .CLK(clknet_leaf_45_clk),
    .Q(\counter6[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0760_ (.D(net213),
    .CLK(clknet_leaf_4_clk),
    .Q(\counter6[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0761_ (.D(net212),
    .CLK(clknet_leaf_4_clk),
    .Q(\counter6[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0762_ (.D(net211),
    .CLK(clknet_leaf_45_clk),
    .Q(\counter6[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0763_ (.D(net210),
    .CLK(clknet_leaf_46_clk),
    .Q(\counter6[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0764_ (.D(net209),
    .CLK(clknet_leaf_46_clk),
    .Q(\counter6[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0765_ (.D(net208),
    .CLK(clknet_leaf_45_clk),
    .Q(\counter6[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0766_ (.D(net207),
    .CLK(clknet_leaf_45_clk),
    .Q(\counter6[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0767_ (.D(net206),
    .CLK(clknet_leaf_47_clk),
    .Q(\counter6[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0768_ (.D(net205),
    .CLK(clknet_leaf_46_clk),
    .Q(\counter6[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0769_ (.D(net204),
    .CLK(clknet_leaf_45_clk),
    .Q(\counter6[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0770_ (.D(net203),
    .CLK(clknet_leaf_47_clk),
    .Q(\counter6[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0771_ (.D(net202),
    .CLK(clknet_leaf_47_clk),
    .Q(\counter6[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0772_ (.D(net201),
    .CLK(clknet_leaf_41_clk),
    .Q(\counter6[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0773_ (.D(net200),
    .CLK(clknet_leaf_41_clk),
    .Q(\counter6[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0774_ (.D(net199),
    .CLK(clknet_leaf_42_clk),
    .Q(\counter6[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0775_ (.D(net198),
    .CLK(clknet_leaf_49_clk),
    .Q(\counter6[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0776_ (.D(net197),
    .CLK(clknet_leaf_49_clk),
    .Q(\counter6[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0777_ (.D(net196),
    .CLK(clknet_leaf_49_clk),
    .Q(\counter6[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0778_ (.D(net195),
    .CLK(clknet_leaf_48_clk),
    .Q(\counter6[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0779_ (.D(net194),
    .CLK(clknet_leaf_48_clk),
    .Q(\counter6[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0780_ (.D(net193),
    .CLK(clknet_leaf_46_clk),
    .Q(\counter6[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0781_ (.D(_0004_),
    .CLK(clknet_leaf_2_clk),
    .Q(net5));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0782_ (.D(_0065_),
    .CLK(clknet_leaf_26_clk),
    .Q(\counter5[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0783_ (.D(_0066_),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\counter5[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0784_ (.D(_0067_),
    .CLK(clknet_leaf_27_clk),
    .Q(\counter5[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0785_ (.D(_0068_),
    .CLK(clknet_leaf_30_clk),
    .Q(\counter5[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0786_ (.D(_0069_),
    .CLK(clknet_leaf_27_clk),
    .Q(\counter5[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0787_ (.D(net192),
    .CLK(clknet_leaf_20_clk),
    .Q(\counter5[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0788_ (.D(net191),
    .CLK(clknet_leaf_20_clk),
    .Q(\counter5[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0789_ (.D(net190),
    .CLK(clknet_leaf_19_clk),
    .Q(\counter5[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0790_ (.D(net189),
    .CLK(clknet_leaf_19_clk),
    .Q(\counter5[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0791_ (.D(net188),
    .CLK(clknet_leaf_19_clk),
    .Q(\counter5[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0792_ (.D(net187),
    .CLK(clknet_leaf_30_clk),
    .Q(\counter5[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0793_ (.D(net186),
    .CLK(clknet_leaf_16_clk),
    .Q(\counter5[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0794_ (.D(net185),
    .CLK(clknet_leaf_22_clk),
    .Q(\counter5[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0795_ (.D(net184),
    .CLK(clknet_leaf_22_clk),
    .Q(\counter5[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0796_ (.D(net183),
    .CLK(clknet_leaf_22_clk),
    .Q(\counter5[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0797_ (.D(net182),
    .CLK(clknet_leaf_18_clk),
    .Q(\counter5[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0798_ (.D(net181),
    .CLK(clknet_leaf_20_clk),
    .Q(\counter5[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0799_ (.D(net180),
    .CLK(clknet_leaf_18_clk),
    .Q(\counter5[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0800_ (.D(net179),
    .CLK(clknet_leaf_19_clk),
    .Q(\counter5[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0801_ (.D(net178),
    .CLK(clknet_leaf_20_clk),
    .Q(\counter5[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0802_ (.D(net177),
    .CLK(clknet_leaf_21_clk),
    .Q(\counter5[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0803_ (.D(net176),
    .CLK(clknet_leaf_30_clk),
    .Q(\counter5[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0804_ (.D(net175),
    .CLK(clknet_leaf_27_clk),
    .Q(\counter5[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0805_ (.D(net174),
    .CLK(clknet_leaf_30_clk),
    .Q(\counter5[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0806_ (.D(net173),
    .CLK(clknet_leaf_30_clk),
    .Q(\counter5[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0807_ (.D(net172),
    .CLK(clknet_leaf_30_clk),
    .Q(\counter5[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0808_ (.D(net171),
    .CLK(clknet_leaf_30_clk),
    .Q(\counter5[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0809_ (.D(net170),
    .CLK(clknet_leaf_20_clk),
    .Q(\counter5[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0810_ (.D(_0003_),
    .CLK(clknet_leaf_40_clk),
    .Q(net4));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0811_ (.D(_0093_),
    .CLK(clknet_leaf_8_clk),
    .Q(\counter4[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0812_ (.D(_0094_),
    .CLK(clknet_leaf_8_clk),
    .Q(\counter4[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0813_ (.D(_0095_),
    .CLK(clknet_leaf_2_clk),
    .Q(\counter4[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0814_ (.D(_0096_),
    .CLK(clknet_leaf_3_clk),
    .Q(\counter4[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0815_ (.D(net169),
    .CLK(clknet_leaf_6_clk),
    .Q(\counter4[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0816_ (.D(net168),
    .CLK(clknet_leaf_18_clk),
    .Q(\counter4[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0817_ (.D(net167),
    .CLK(clknet_leaf_5_clk),
    .Q(\counter4[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0818_ (.D(net166),
    .CLK(clknet_leaf_19_clk),
    .Q(\counter4[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0819_ (.D(net165),
    .CLK(clknet_leaf_5_clk),
    .Q(\counter4[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0820_ (.D(net164),
    .CLK(clknet_leaf_6_clk),
    .Q(\counter4[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0821_ (.D(net163),
    .CLK(clknet_leaf_5_clk),
    .Q(\counter4[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0822_ (.D(net162),
    .CLK(clknet_leaf_5_clk),
    .Q(\counter4[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0823_ (.D(net161),
    .CLK(clknet_leaf_6_clk),
    .Q(\counter4[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0824_ (.D(net160),
    .CLK(clknet_leaf_6_clk),
    .Q(\counter4[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0825_ (.D(net159),
    .CLK(clknet_leaf_6_clk),
    .Q(\counter4[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0826_ (.D(net158),
    .CLK(clknet_leaf_6_clk),
    .Q(\counter4[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0827_ (.D(net157),
    .CLK(clknet_leaf_4_clk),
    .Q(\counter4[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0828_ (.D(net156),
    .CLK(clknet_leaf_4_clk),
    .Q(\counter4[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0829_ (.D(net155),
    .CLK(clknet_leaf_4_clk),
    .Q(\counter4[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0830_ (.D(net154),
    .CLK(clknet_leaf_4_clk),
    .Q(\counter4[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0831_ (.D(net153),
    .CLK(clknet_leaf_8_clk),
    .Q(\counter4[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0832_ (.D(net152),
    .CLK(clknet_leaf_3_clk),
    .Q(\counter4[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0833_ (.D(net151),
    .CLK(clknet_leaf_3_clk),
    .Q(\counter4[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0834_ (.D(net150),
    .CLK(clknet_leaf_3_clk),
    .Q(\counter4[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0835_ (.D(net149),
    .CLK(clknet_leaf_7_clk),
    .Q(\counter4[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0836_ (.D(net148),
    .CLK(clknet_leaf_8_clk),
    .Q(\counter4[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0837_ (.D(net147),
    .CLK(clknet_leaf_7_clk),
    .Q(\counter4[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0838_ (.D(net146),
    .CLK(clknet_leaf_7_clk),
    .Q(\counter4[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0839_ (.D(_0002_),
    .CLK(clknet_leaf_25_clk),
    .Q(net3));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0840_ (.D(_0121_),
    .CLK(clknet_leaf_42_clk),
    .Q(\counter3[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0841_ (.D(_0122_),
    .CLK(clknet_leaf_40_clk),
    .Q(\counter3[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0842_ (.D(_0123_),
    .CLK(clknet_leaf_40_clk),
    .Q(\counter3[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0843_ (.D(net145),
    .CLK(clknet_leaf_42_clk),
    .Q(\counter3[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0844_ (.D(net144),
    .CLK(clknet_leaf_42_clk),
    .Q(\counter3[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0845_ (.D(net143),
    .CLK(clknet_leaf_43_clk),
    .Q(\counter3[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0846_ (.D(net142),
    .CLK(clknet_leaf_43_clk),
    .Q(\counter3[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0847_ (.D(net141),
    .CLK(clknet_leaf_33_clk),
    .Q(\counter3[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0848_ (.D(net140),
    .CLK(clknet_leaf_43_clk),
    .Q(\counter3[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0849_ (.D(net139),
    .CLK(clknet_leaf_41_clk),
    .Q(\counter3[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0850_ (.D(net138),
    .CLK(clknet_leaf_45_clk),
    .Q(\counter3[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0851_ (.D(net137),
    .CLK(clknet_leaf_43_clk),
    .Q(\counter3[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0852_ (.D(net136),
    .CLK(clknet_leaf_41_clk),
    .Q(\counter3[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0853_ (.D(net135),
    .CLK(clknet_leaf_43_clk),
    .Q(\counter3[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0854_ (.D(net134),
    .CLK(clknet_leaf_32_clk),
    .Q(\counter3[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0855_ (.D(net133),
    .CLK(clknet_leaf_43_clk),
    .Q(\counter3[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0856_ (.D(net132),
    .CLK(clknet_leaf_32_clk),
    .Q(\counter3[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0857_ (.D(net131),
    .CLK(clknet_leaf_5_clk),
    .Q(\counter3[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0858_ (.D(net130),
    .CLK(clknet_leaf_19_clk),
    .Q(\counter3[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0859_ (.D(net129),
    .CLK(clknet_leaf_5_clk),
    .Q(\counter3[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0860_ (.D(net128),
    .CLK(clknet_leaf_19_clk),
    .Q(\counter3[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0861_ (.D(net127),
    .CLK(clknet_leaf_5_clk),
    .Q(\counter3[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0862_ (.D(net126),
    .CLK(clknet_leaf_44_clk),
    .Q(\counter3[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0863_ (.D(net125),
    .CLK(clknet_leaf_44_clk),
    .Q(\counter3[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0864_ (.D(net124),
    .CLK(clknet_leaf_44_clk),
    .Q(\counter3[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0865_ (.D(net123),
    .CLK(clknet_leaf_43_clk),
    .Q(\counter3[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0866_ (.D(net122),
    .CLK(clknet_leaf_44_clk),
    .Q(\counter3[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0867_ (.D(net121),
    .CLK(clknet_leaf_42_clk),
    .Q(\counter3[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0868_ (.D(_0001_),
    .CLK(clknet_leaf_38_clk),
    .Q(net1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0869_ (.D(_0149_),
    .CLK(clknet_leaf_25_clk),
    .Q(\counter2[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0870_ (.D(_0150_),
    .CLK(clknet_leaf_25_clk),
    .Q(\counter2[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0871_ (.D(net120),
    .CLK(clknet_leaf_25_clk),
    .Q(\counter2[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0872_ (.D(net119),
    .CLK(clknet_leaf_25_clk),
    .Q(\counter2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0873_ (.D(net118),
    .CLK(clknet_leaf_25_clk),
    .Q(\counter2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0874_ (.D(net117),
    .CLK(clknet_leaf_25_clk),
    .Q(\counter2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0875_ (.D(net116),
    .CLK(clknet_leaf_26_clk),
    .Q(\counter2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0876_ (.D(net115),
    .CLK(clknet_leaf_26_clk),
    .Q(\counter2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0877_ (.D(net114),
    .CLK(clknet_leaf_25_clk),
    .Q(\counter2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0878_ (.D(net113),
    .CLK(clknet_leaf_26_clk),
    .Q(\counter2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0879_ (.D(net112),
    .CLK(clknet_leaf_24_clk),
    .Q(\counter2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0880_ (.D(net111),
    .CLK(clknet_leaf_24_clk),
    .Q(\counter2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0881_ (.D(net110),
    .CLK(clknet_leaf_26_clk),
    .Q(\counter2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0882_ (.D(net109),
    .CLK(clknet_leaf_25_clk),
    .Q(\counter2[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0883_ (.D(net108),
    .CLK(clknet_leaf_21_clk),
    .Q(\counter2[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0884_ (.D(net107),
    .CLK(clknet_leaf_21_clk),
    .Q(\counter2[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0885_ (.D(net106),
    .CLK(clknet_leaf_21_clk),
    .Q(\counter2[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0886_ (.D(net105),
    .CLK(clknet_leaf_24_clk),
    .Q(\counter2[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0887_ (.D(net104),
    .CLK(clknet_leaf_24_clk),
    .Q(\counter2[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0888_ (.D(net103),
    .CLK(clknet_leaf_22_clk),
    .Q(\counter2[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0889_ (.D(net102),
    .CLK(clknet_leaf_24_clk),
    .Q(\counter2[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0890_ (.D(net101),
    .CLK(clknet_leaf_23_clk),
    .Q(\counter2[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0891_ (.D(net100),
    .CLK(clknet_leaf_23_clk),
    .Q(\counter2[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0892_ (.D(net99),
    .CLK(clknet_leaf_23_clk),
    .Q(\counter2[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0893_ (.D(net98),
    .CLK(clknet_leaf_23_clk),
    .Q(\counter2[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0894_ (.D(net97),
    .CLK(clknet_leaf_23_clk),
    .Q(\counter2[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0895_ (.D(net96),
    .CLK(clknet_leaf_23_clk),
    .Q(\counter2[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0896_ (.D(net95),
    .CLK(clknet_leaf_23_clk),
    .Q(\counter2[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0897_ (.D(_0000_),
    .CLK(clknet_leaf_50_clk),
    .Q(net2));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0898_ (.D(_0177_),
    .CLK(clknet_leaf_37_clk),
    .Q(\counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0899_ (.D(net94),
    .CLK(clknet_leaf_38_clk),
    .Q(\counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0900_ (.D(net93),
    .CLK(clknet_leaf_39_clk),
    .Q(\counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0901_ (.D(net92),
    .CLK(clknet_leaf_39_clk),
    .Q(\counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0902_ (.D(net91),
    .CLK(clknet_leaf_36_clk),
    .Q(\counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0903_ (.D(net90),
    .CLK(clknet_leaf_40_clk),
    .Q(\counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0904_ (.D(net89),
    .CLK(clknet_leaf_40_clk),
    .Q(\counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0905_ (.D(net88),
    .CLK(clknet_leaf_40_clk),
    .Q(\counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0906_ (.D(net87),
    .CLK(clknet_leaf_38_clk),
    .Q(\counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0907_ (.D(net86),
    .CLK(clknet_leaf_36_clk),
    .Q(\counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0908_ (.D(net85),
    .CLK(clknet_leaf_42_clk),
    .Q(\counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0909_ (.D(net84),
    .CLK(clknet_leaf_33_clk),
    .Q(\counter[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0910_ (.D(net83),
    .CLK(clknet_leaf_36_clk),
    .Q(\counter[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0911_ (.D(net82),
    .CLK(clknet_leaf_36_clk),
    .Q(\counter[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0912_ (.D(net81),
    .CLK(clknet_leaf_36_clk),
    .Q(\counter[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0913_ (.D(net80),
    .CLK(clknet_leaf_36_clk),
    .Q(\counter[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0914_ (.D(net79),
    .CLK(clknet_leaf_37_clk),
    .Q(\counter[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0915_ (.D(net78),
    .CLK(clknet_leaf_36_clk),
    .Q(\counter[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0916_ (.D(net77),
    .CLK(clknet_leaf_36_clk),
    .Q(\counter[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0917_ (.D(net76),
    .CLK(clknet_leaf_35_clk),
    .Q(\counter[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0918_ (.D(net75),
    .CLK(clknet_leaf_35_clk),
    .Q(\counter[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0919_ (.D(net74),
    .CLK(clknet_leaf_38_clk),
    .Q(\counter[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0920_ (.D(net73),
    .CLK(clknet_leaf_38_clk),
    .Q(\counter[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0921_ (.D(net72),
    .CLK(clknet_leaf_38_clk),
    .Q(\counter[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0922_ (.D(net71),
    .CLK(clknet_leaf_37_clk),
    .Q(\counter[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0923_ (.D(net70),
    .CLK(clknet_leaf_38_clk),
    .Q(\counter[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0924_ (.D(net69),
    .CLK(clknet_leaf_37_clk),
    .Q(\counter[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0925_ (.D(net68),
    .CLK(clknet_leaf_39_clk),
    .Q(\counter[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0926_ (.D(_0009_),
    .CLK(clknet_leaf_34_clk),
    .Q(net10));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0927_ (.D(_0205_),
    .CLK(clknet_leaf_50_clk),
    .Q(\counter10[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0928_ (.D(_0206_),
    .CLK(clknet_leaf_0_clk),
    .Q(\counter10[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0929_ (.D(_0207_),
    .CLK(clknet_leaf_0_clk),
    .Q(\counter10[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0930_ (.D(_0208_),
    .CLK(clknet_leaf_50_clk),
    .Q(\counter10[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0931_ (.D(_0209_),
    .CLK(clknet_leaf_50_clk),
    .Q(\counter10[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0932_ (.D(_0210_),
    .CLK(clknet_leaf_49_clk),
    .Q(\counter10[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0933_ (.D(_0211_),
    .CLK(clknet_leaf_49_clk),
    .Q(\counter10[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0934_ (.D(_0212_),
    .CLK(clknet_leaf_49_clk),
    .Q(\counter10[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0935_ (.D(_0213_),
    .CLK(clknet_leaf_1_clk),
    .Q(\counter10[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0936_ (.D(_0214_),
    .CLK(clknet_leaf_0_clk),
    .Q(\counter10[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0937_ (.D(net67),
    .CLK(clknet_leaf_1_clk),
    .Q(\counter10[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0938_ (.D(net66),
    .CLK(clknet_leaf_1_clk),
    .Q(\counter10[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0939_ (.D(net65),
    .CLK(clknet_leaf_1_clk),
    .Q(\counter10[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0940_ (.D(net64),
    .CLK(clknet_leaf_49_clk),
    .Q(\counter10[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0941_ (.D(net63),
    .CLK(clknet_leaf_2_clk),
    .Q(\counter10[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0942_ (.D(net62),
    .CLK(clknet_leaf_3_clk),
    .Q(\counter10[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0943_ (.D(net61),
    .CLK(clknet_leaf_1_clk),
    .Q(\counter10[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0944_ (.D(net60),
    .CLK(clknet_leaf_3_clk),
    .Q(\counter10[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0945_ (.D(net59),
    .CLK(clknet_leaf_3_clk),
    .Q(\counter10[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0946_ (.D(net58),
    .CLK(clknet_leaf_4_clk),
    .Q(\counter10[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0947_ (.D(net57),
    .CLK(clknet_leaf_3_clk),
    .Q(\counter10[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0948_ (.D(net56),
    .CLK(clknet_leaf_4_clk),
    .Q(\counter10[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0949_ (.D(net55),
    .CLK(clknet_leaf_2_clk),
    .Q(\counter10[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0950_ (.D(net54),
    .CLK(clknet_leaf_2_clk),
    .Q(\counter10[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0951_ (.D(net53),
    .CLK(clknet_leaf_2_clk),
    .Q(\counter10[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0952_ (.D(net52),
    .CLK(clknet_leaf_2_clk),
    .Q(\counter10[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0953_ (.D(net51),
    .CLK(clknet_leaf_1_clk),
    .Q(\counter10[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0954_ (.D(net50),
    .CLK(clknet_leaf_1_clk),
    .Q(\counter10[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0955_ (.D(_0008_),
    .CLK(clknet_leaf_15_clk),
    .Q(net9));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0956_ (.D(_0233_),
    .CLK(clknet_leaf_33_clk),
    .Q(\counter9[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0957_ (.D(_0234_),
    .CLK(clknet_leaf_33_clk),
    .Q(\counter9[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0958_ (.D(_0235_),
    .CLK(clknet_leaf_33_clk),
    .Q(\counter9[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0959_ (.D(_0236_),
    .CLK(clknet_leaf_36_clk),
    .Q(\counter9[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0960_ (.D(_0237_),
    .CLK(clknet_leaf_36_clk),
    .Q(\counter9[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0961_ (.D(_0238_),
    .CLK(clknet_leaf_35_clk),
    .Q(\counter9[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0962_ (.D(_0239_),
    .CLK(clknet_leaf_35_clk),
    .Q(\counter9[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0963_ (.D(_0240_),
    .CLK(clknet_leaf_34_clk),
    .Q(\counter9[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0964_ (.D(_0241_),
    .CLK(clknet_leaf_34_clk),
    .Q(\counter9[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0965_ (.D(net49),
    .CLK(clknet_leaf_33_clk),
    .Q(\counter9[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0966_ (.D(net48),
    .CLK(clknet_leaf_33_clk),
    .Q(\counter9[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0967_ (.D(net47),
    .CLK(clknet_leaf_31_clk),
    .Q(\counter9[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0968_ (.D(net46),
    .CLK(clknet_leaf_32_clk),
    .Q(\counter9[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0969_ (.D(net45),
    .CLK(clknet_leaf_31_clk),
    .Q(\counter9[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0970_ (.D(net44),
    .CLK(clknet_leaf_31_clk),
    .Q(\counter9[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0971_ (.D(net43),
    .CLK(clknet_leaf_32_clk),
    .Q(\counter9[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0972_ (.D(net42),
    .CLK(clknet_leaf_32_clk),
    .Q(\counter9[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0973_ (.D(net41),
    .CLK(clknet_leaf_32_clk),
    .Q(\counter9[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0974_ (.D(net40),
    .CLK(clknet_leaf_33_clk),
    .Q(\counter9[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0975_ (.D(net39),
    .CLK(clknet_leaf_30_clk),
    .Q(\counter9[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0976_ (.D(net38),
    .CLK(clknet_leaf_31_clk),
    .Q(\counter9[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0977_ (.D(net37),
    .CLK(clknet_leaf_30_clk),
    .Q(\counter9[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0978_ (.D(net36),
    .CLK(clknet_leaf_34_clk),
    .Q(\counter9[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0979_ (.D(net35),
    .CLK(clknet_leaf_30_clk),
    .Q(\counter9[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0980_ (.D(net34),
    .CLK(clknet_leaf_29_clk),
    .Q(\counter9[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0981_ (.D(net33),
    .CLK(clknet_leaf_29_clk),
    .Q(\counter9[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0982_ (.D(net32),
    .CLK(clknet_leaf_29_clk),
    .Q(\counter9[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0983_ (.D(net31),
    .CLK(clknet_leaf_33_clk),
    .Q(\counter9[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0984_ (.D(_0007_),
    .CLK(clknet_leaf_12_clk),
    .Q(net8));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0985_ (.D(_0261_),
    .CLK(clknet_leaf_15_clk),
    .Q(\counter8[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0986_ (.D(_0262_),
    .CLK(clknet_leaf_15_clk),
    .Q(\counter8[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0987_ (.D(_0263_),
    .CLK(clknet_leaf_22_clk),
    .Q(\counter8[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0988_ (.D(_0264_),
    .CLK(clknet_leaf_15_clk),
    .Q(\counter8[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0989_ (.D(_0265_),
    .CLK(clknet_leaf_16_clk),
    .Q(\counter8[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0990_ (.D(_0266_),
    .CLK(clknet_leaf_17_clk),
    .Q(\counter8[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0991_ (.D(_0267_),
    .CLK(clknet_leaf_15_clk),
    .Q(\counter8[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0992_ (.D(_0268_),
    .CLK(clknet_leaf_15_clk),
    .Q(\counter8[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0993_ (.D(net30),
    .CLK(clknet_leaf_17_clk),
    .Q(\counter8[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0994_ (.D(net29),
    .CLK(clknet_leaf_17_clk),
    .Q(\counter8[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0995_ (.D(net28),
    .CLK(clknet_leaf_17_clk),
    .Q(\counter8[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0996_ (.D(net27),
    .CLK(clknet_leaf_17_clk),
    .Q(\counter8[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0997_ (.D(net26),
    .CLK(clknet_leaf_18_clk),
    .Q(\counter8[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0998_ (.D(net25),
    .CLK(clknet_leaf_18_clk),
    .Q(\counter8[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _0999_ (.D(net24),
    .CLK(clknet_leaf_16_clk),
    .Q(\counter8[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1000_ (.D(net23),
    .CLK(clknet_leaf_18_clk),
    .Q(\counter8[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1001_ (.D(net22),
    .CLK(clknet_leaf_7_clk),
    .Q(\counter8[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1002_ (.D(net21),
    .CLK(clknet_leaf_6_clk),
    .Q(\counter8[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1003_ (.D(net20),
    .CLK(clknet_leaf_17_clk),
    .Q(\counter8[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1004_ (.D(net19),
    .CLK(clknet_leaf_6_clk),
    .Q(\counter8[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1005_ (.D(net18),
    .CLK(clknet_leaf_14_clk),
    .Q(\counter8[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1006_ (.D(net17),
    .CLK(clknet_leaf_14_clk),
    .Q(\counter8[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1007_ (.D(net16),
    .CLK(clknet_leaf_13_clk),
    .Q(\counter8[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1008_ (.D(net15),
    .CLK(clknet_leaf_14_clk),
    .Q(\counter8[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1009_ (.D(net14),
    .CLK(clknet_leaf_14_clk),
    .Q(\counter8[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1010_ (.D(net13),
    .CLK(clknet_leaf_13_clk),
    .Q(\counter8[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1011_ (.D(net12),
    .CLK(clknet_leaf_14_clk),
    .Q(\counter8[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1012_ (.D(net11),
    .CLK(clknet_leaf_14_clk),
    .Q(\counter8[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1013_ (.D(_0006_),
    .CLK(clknet_leaf_48_clk),
    .Q(net7));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1014_ (.D(_0289_),
    .CLK(clknet_leaf_13_clk),
    .Q(\counter7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1011__12 (.ZN(net12));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1010__13 (.ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1009__14 (.ZN(net14));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1008__15 (.ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1007__16 (.ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1006__17 (.ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1005__18 (.ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1004__19 (.ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1003__20 (.ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1002__21 (.ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1001__22 (.ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1000__23 (.ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0999__24 (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0998__25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0997__26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0996__27 (.ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0995__28 (.ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0994__29 (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0993__30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0983__31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0982__32 (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0981__33 (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0980__34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0979__35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0978__36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0977__37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0976__38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0975__39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0974__40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0973__41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0972__42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0971__43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0970__44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0969__45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0968__46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0967__47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0966__48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0965__49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0954__50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0953__51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0952__52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0951__53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0950__54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0949__55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0948__56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0947__57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0946__58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0945__59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0944__60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0943__61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0942__62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0941__63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0940__64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0939__65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0938__66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0937__67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0925__68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0924__69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0923__70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0922__71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0921__72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0920__73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0919__74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0918__75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0917__76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0916__77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0915__78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0914__79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0913__80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0912__81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0911__82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0910__83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0909__84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0908__85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0907__86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0906__87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0905__88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0904__89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0903__90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0902__91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0901__92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0900__93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0899__94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0896__95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0895__96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0894__97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0893__98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0892__99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0891__100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0890__101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0889__102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0888__103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0887__104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0886__105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0885__106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0884__107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0883__108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0882__109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0881__110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0880__111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0879__112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0878__113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0877__114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0876__115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0875__116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0874__117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0873__118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0872__119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0871__120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0867__121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0866__122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0865__123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0864__124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0863__125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0862__126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0861__127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0860__128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0859__129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0858__130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0857__131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0856__132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0855__133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0854__134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0853__135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0852__136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0851__137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0850__138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0849__139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0848__140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0847__141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0846__142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0845__143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0844__144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0843__145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0838__146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0837__147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0836__148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0835__149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0834__150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0833__151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0832__152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0831__153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0830__154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0829__155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0828__156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0827__157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0826__158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0825__159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0824__160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0823__161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0822__162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0821__163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0820__164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0819__165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0818__166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0817__167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0816__168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0815__169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0809__170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0808__171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0807__172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0806__173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0805__174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0804__175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0803__176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0802__177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0801__178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0800__179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0799__180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0798__181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0797__182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0796__183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0795__184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0794__185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0793__186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0792__187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0791__188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0790__189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0789__190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0788__191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0787__192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0780__193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0779__194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0778__195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0777__196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0776__197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0775__198 (.ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0774__199 (.ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0773__200 (.ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0772__201 (.ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0771__202 (.ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0770__203 (.ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0769__204 (.ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0768__205 (.ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0767__206 (.ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0766__207 (.ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0765__208 (.ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0764__209 (.ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0763__210 (.ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0762__211 (.ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0761__212 (.ZN(net212));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0760__213 (.ZN(net213));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0759__214 (.ZN(net214));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0751__215 (.ZN(net215));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0750__216 (.ZN(net216));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0749__217 (.ZN(net217));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0748__218 (.ZN(net218));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0747__219 (.ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0746__220 (.ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0745__221 (.ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0744__222 (.ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0743__223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0742__224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0741__225 (.ZN(net225));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0740__226 (.ZN(net226));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0739__227 (.ZN(net227));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0738__228 (.ZN(net228));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0737__229 (.ZN(net229));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0736__230 (.ZN(net230));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0735__231 (.ZN(net231));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0734__232 (.ZN(net232));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0733__233 (.ZN(net233));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0732__234 (.ZN(net234));
 gf180mcu_fd_sc_mcu7t5v0__tiel _0731__235 (.ZN(net235));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output1 (.I(net1),
    .Z(cout1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output2 (.I(net2),
    .Z(cout10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output3 (.I(net3),
    .Z(cout2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output4 (.I(net4),
    .Z(cout3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output5 (.I(net5),
    .Z(cout4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output6 (.I(net6),
    .Z(cout5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(cout6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output8 (.I(net8),
    .Z(cout7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output9 (.I(net9),
    .Z(cout8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output10 (.I(net10),
    .Z(cout9));
 gf180mcu_fd_sc_mcu7t5v0__tiel _1012__11 (.ZN(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_16_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_29_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clk (.I(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clk (.I(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0752__D (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0719__A2 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0714__A2 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0711__A2 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0705__I (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0723__B (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0716__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0708__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0706__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0493__A2 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0503__A4 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0636__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0633__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0631__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0504__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0630__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0513__I (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0589__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0586__A1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0543__A2 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0697__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0676__B (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0561__A3 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0671__B2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0650__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0648__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0572__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0607__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0600__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0598__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0595__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0666__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0663__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0656__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0644__A3 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0665__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0660__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0650__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0648__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output8_I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0953__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0954__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0943__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0938__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0939__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0935__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0937__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0813__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0950__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0941__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0949__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0781__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0951__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0952__CLK (.I(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0947__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0942__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0833__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0945__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0834__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0832__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0944__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0814__CLK (.I(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0828__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0830__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0829__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0760__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0761__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0827__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0948__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0946__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0817__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0857__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0859__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0822__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0861__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0819__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0821__CLK (.I(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1002__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1004__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0824__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0823__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0826__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0825__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0820__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0815__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0835__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0838__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0837__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0743__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0738__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0737__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1001__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0744__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0812__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0836__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0811__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0831__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0740__CLK (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0746__CLK (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0742__CLK (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0747__CLK (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0741__CLK (.I(clknet_leaf_9_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0745__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0748__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0735__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0736__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0739__CLK (.I(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0731__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0728__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0749__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0750__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0732__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0751__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0734__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1010__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1007__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1014__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0727__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1005__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1006__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0725__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1008__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0726__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1009__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1011__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0733__CLK (.I(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0988__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0985__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0991__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0986__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0955__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0992__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0995__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0993__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0994__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0996__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0990__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0816__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0799__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0797__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0997__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1000__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0998__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0800__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0789__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0791__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0790__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0858__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0860__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0818__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0801__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0788__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0787__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0809__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0798__CLK (.I(clknet_leaf_20_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0987__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0888__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0794__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0796__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0795__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0896__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0895__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0890__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0893__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0892__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0894__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0891__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0879__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0880__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0886__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0887__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0889__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0877__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0752__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0874__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0872__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0873__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0870__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0839__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0882__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0869__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0871__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0876__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0881__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0875__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0782__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0878__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0975__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0977__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0807__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0806__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0792__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0805__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0803__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0808__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0979__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0785__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0967__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0970__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0969__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0976__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0957__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0909__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0847__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0958__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0966__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0965__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0983__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0956__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0974__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0926__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0963__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0964__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0978__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0918__CLK (.I(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0917__CLK (.I(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0961__CLK (.I(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0962__CLK (.I(clknet_leaf_35_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0902__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0912__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0911__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0907__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0910__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0916__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0915__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0959__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0960__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0913__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0922__CLK (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0924__CLK (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0914__CLK (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0898__CLK (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0899__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0906__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0920__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0921__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0919__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0923__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0868__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0842__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0810__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0905__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0904__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0903__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0841__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0852__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0849__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0773__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0772__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0754__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0908__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0844__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0774__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0840__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0867__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0843__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0855__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0848__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0853__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0865__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0851__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0846__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0845__CLK (.I(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0765__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0759__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0762__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0766__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0769__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0850__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0780__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0768__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0764__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0763__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0779__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0757__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0778__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0758__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1013__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0756__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0753__CLK (.I(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0932__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0933__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0934__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0776__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0940__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0775__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0777__CLK (.I(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clk_I (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0783__CLK (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clk_I (.I(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_508 ();
endmodule

