* NGSPICE file created from divider.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

.subckt divider clk cout1 cout10 cout2 cout3 cout4 cout5 cout6 cout7 cout8 cout9 vdd
+ vss
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0949__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0965__49 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0985_ _0261_ clknet_leaf_15_clk counter8\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0650__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0770_ net203 clknet_leaf_47_clk counter6\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0794__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0968_ net46 clknet_leaf_32_clk counter9\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0899_ net94 clknet_leaf_38_clk counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0952__52 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_55_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0822_ net162 clknet_leaf_5_clk counter4\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0684_ _0463_ _0464_ _0465_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0753_ _0037_ clknet_leaf_48_clk counter6\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_37_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0656__I _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0832__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0805_ net174 clknet_leaf_30_clk counter5\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0736_ net230 clknet_leaf_10_clk counter7\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0598_ _0410_ _0409_ _0411_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0667_ counter10\[7\] _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0855__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0521_ _0344_ _0345_ _0346_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1010__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1004_ net19 clknet_leaf_6_clk counter8\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0728__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0878__CLK clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0719_ _0302_ _0294_ _0303_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput7 net7 cout6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0837__147 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0504_ counter3\[2\] _0332_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0708__A1 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0984_ _0007_ clknet_leaf_12_clk net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0916__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0827__157 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0939__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0967_ net47 clknet_leaf_31_clk counter9\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0898_ _0177_ clknet_leaf_37_clk counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0752_ _0005_ clknet_leaf_25_clk net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0821_ net163 clknet_leaf_5_clk counter4\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0683_ counter9\[1\] _0456_ counter9\[2\] _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__0761__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0817__167 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0735_ net231 clknet_leaf_10_clk counter7\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0804_ net175 clknet_leaf_27_clk counter5\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0597_ counter6\[1\] counter6\[0\] _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0666_ counter10\[6\] _0436_ _0437_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0907__86 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_49_clk clknet_2_0__leaf_clk clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0798__181 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0520_ counter5\[6\] counter5\[5\] counter5\[27\] _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_21_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1003_ net20 clknet_leaf_17_clk counter8\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0904__89 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_19_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_36_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0718_ counter8\[4\] _0299_ counter8\[5\] _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0649_ counter10\[1\] _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0977__37 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xoutput8 net8 cout7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput10 net10 cout9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__0822__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0671__B2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0503_ _0324_ _0325_ _0326_ _0331_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_50_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0788__191 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0845__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0795__184 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_45_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0995__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1000__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0983_ net31 clknet_leaf_33_clk counter9\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0868__CLK clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0966_ net48 clknet_leaf_33_clk counter9\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0897_ _0000_ clknet_leaf_50_clk net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0792__187 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_28_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0833__151 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0751_ net215 clknet_leaf_11_clk counter7\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0820_ net164 clknet_leaf_6_clk counter4\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0682_ _0460_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0906__CLK clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1009__14 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_52_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0748__218 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0949_ net55 clknet_leaf_2_clk counter10\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1006__17 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0734_ net232 clknet_leaf_13_clk counter7\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0803_ net176 clknet_leaf_30_clk counter5\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0665_ _0448_ _0440_ _0452_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0823__161 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0596_ counter6\[1\] counter6\[0\] _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_37_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0830__154 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0751__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0738__228 net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1002_ net21 clknet_leaf_6_clk counter8\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0717_ counter8\[4\] counter8\[5\] _0299_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_0648_ _0393_ _0440_ _0441_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0579_ _0394_ _0398_ _0399_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_57_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0903__90 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_25_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0774__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput9 net9 cout8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0502_ _0327_ _0328_ _0329_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__0797__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0820__164 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0900__93 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_30_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_20_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0973__41 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_clkbuf_leaf_35_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0982_ net32 clknet_leaf_29_clk counter9\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0812__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0962__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0970__44 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_61_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0835__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0896_ net95 clknet_leaf_23_clk counter2\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0985__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0965_ net49 clknet_leaf_33_clk counter9\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0858__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_2_2__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0750_ net216 clknet_leaf_11_clk counter7\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0681_ counter9\[2\] counter9\[1\] _0456_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_6_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0919__74 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1013__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0948_ net56 clknet_leaf_4_clk counter10\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0879_ net112 clknet_leaf_24_clk counter2\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0916__77 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0802_ net177 clknet_leaf_21_clk counter5\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0998__25 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0733_ net233 clknet_leaf_14_clk counter7\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0664_ counter10\[6\] _0451_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_0595_ counter6\[0\] _0409_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0995__28 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1001_ net22 clknet_leaf_7_clk counter8\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0578_ counter7\[0\] counter7\[1\] _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0716_ _0295_ _0301_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1002__21 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0647_ counter10\[0\] _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0919__CLK clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_9_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0744__222 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0501_ counter3\[16\] counter3\[15\] counter3\[14\] counter3\[13\] _0330_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0751__215 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0741__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0891__CLK clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0981_ net33 clknet_leaf_29_clk counter9\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0644__A3 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0764__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_clk clknet_2_3__leaf_clk clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0734__232 net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__0787__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0741__225 net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_12_clk clknet_2_1__leaf_clk clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0964_ _0241_ clknet_leaf_34_clk counter9\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0895_ net96 clknet_leaf_23_clk counter2\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_34_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_49_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0680_ _0461_ _0462_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0952__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0947_ net57 clknet_leaf_3_clk counter10\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0878_ net113 clknet_leaf_26_clk counter2\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0731__235 net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0825__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0975__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0801_ net178 clknet_leaf_20_clk counter5\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0732_ net234 clknet_leaf_11_clk counter7\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0663_ _0436_ _0437_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0594_ _0352_ _0355_ _0358_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_25_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0848__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0998__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1003__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1000_ net23 clknet_leaf_18_clk counter8\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0912__81 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_19_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0715_ counter8\[4\] _0299_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0577_ _0397_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0646_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0500_ counter3\[20\] counter3\[19\] counter3\[18\] counter3\[17\] _0329_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0982__32 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_30_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0629_ counter4\[3\] _0427_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0980_ net34 clknet_leaf_29_clk counter9\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0909__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0866__122 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_8_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0894_ net97 clknet_leaf_23_clk counter2\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0731__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0963_ _0240_ clknet_leaf_34_clk counter9\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0881__CLK clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0754__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0856__132 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0877_ net114 clknet_leaf_25_clk counter2\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0863__125 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0946_ net58 clknet_leaf_4_clk counter10\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0925__68 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0777__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0731_ net235 clknet_leaf_11_clk counter7\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0800_ net179 clknet_leaf_19_clk counter5\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_33_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0662_ _0447_ _0437_ _0439_ _0448_ _0450_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_0593_ counter6\[5\] counter6\[4\] _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_48_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0929_ _0207_ clknet_leaf_0_clk counter10\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0846__142 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1011__12 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0942__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0853__135 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0714_ _0299_ _0294_ _0300_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0860__128 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0645_ _0435_ _0438_ _0391_ _0387_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_0576_ _0361_ _0364_ _0366_ _0396_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0665__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0815__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0965__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0838__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0988__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0628_ counter4\[3\] _0427_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0559_ counter9\[18\] counter9\[17\] counter9\[16\] counter9\[15\] _0382_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0843__145 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0850__138 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0893_ net98 clknet_leaf_23_clk counter2\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0962_ _0239_ clknet_leaf_35_clk counter9\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0876_ net115 clknet_leaf_26_clk counter2\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_7_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0945_ net59 clknet_leaf_3_clk counter10\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0871__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0730_ _0015_ clknet_leaf_12_clk counter7\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0661_ counter10\[4\] _0447_ counter10\[5\] _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0592_ counter6\[1\] counter6\[0\] counter6\[2\] counter6\[3\] _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0744__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0859_ net129 clknet_leaf_5_clk counter3\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0928_ _0206_ clknet_leaf_0_clk counter10\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0894__CLK clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0921__72 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0713_ counter8\[3\] _0297_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0644_ counter10\[7\] counter10\[6\] _0436_ _0437_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_0575_ counter7\[6\] counter7\[5\] counter7\[4\] _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_38_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_32_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_47_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_42_clk clknet_2_2__leaf_clk clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0558_ counter9\[14\] counter9\[13\] counter9\[12\] counter9\[11\] _0381_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_0627_ _0341_ _0427_ _0428_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0489_ counter2\[25\] counter2\[24\] counter2\[23\] counter2\[22\] _0319_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_38_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_33_clk clknet_2_2__leaf_clk clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__0932__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_24_clk clknet_2_3__leaf_clk clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0805__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0955__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_15_clk clknet_2_1__leaf_clk clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_50_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0828__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0978__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0778__195 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0889__102 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0961_ _0238_ clknet_leaf_35_clk counter9\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0892_ net99 clknet_leaf_23_clk counter2\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_4_clk clknet_2_0__leaf_clk clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0937__67 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_55_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1006__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0676__B _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0944_ net60 clknet_leaf_3_clk counter10\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0875_ net116 clknet_leaf_26_clk counter2\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0752__D _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0879__112 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_46_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0775__198 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_19_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0886__105 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_42_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0591_ _0398_ _0406_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0660_ _0448_ _0440_ _0449_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0927_ _0205_ clknet_leaf_50_clk counter10\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0789_ net190 clknet_leaf_19_clk counter5\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0858_ net130 clknet_leaf_19_clk counter3\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_6_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0574_ counter7\[0\] counter7\[3\] counter7\[2\] counter7\[1\] _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_0712_ _0292_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0643_ counter10\[5\] counter10\[4\] _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0876__115 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0861__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0883__108 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_12_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0734__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_clk clk clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0626_ counter4\[2\] _0425_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0557_ counter9\[10\] counter9\[9\] counter9\[27\] _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0488_ counter2\[1\] counter2\[0\] counter2\[27\] counter2\[26\] _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0894__97 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0757__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0873__118 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0609_ counter5\[3\] _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_31_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_46_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0960_ _0237_ clknet_leaf_36_clk counter9\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0891_ net100 clknet_leaf_23_clk counter2\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0922__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0945__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0874_ net117 clknet_leaf_25_clk counter2\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0943_ net61 clknet_leaf_1_clk counter10\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0818__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0809__170 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_59_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0590_ counter7\[5\] _0402_ counter7\[6\] _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0857_ net131 clknet_leaf_5_clk counter3\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0926_ _0009_ clknet_leaf_34_clk net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0788_ net191 clknet_leaf_20_clk counter5\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0790__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0711_ _0297_ _0294_ _0298_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0573_ counter7\[0\] counter7\[1\] _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_0642_ counter10\[1\] counter10\[0\] counter10\[3\] counter10\[2\] _0436_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0586__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0909_ net84 clknet_leaf_33_clk counter\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0806__173 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0625_ counter4\[2\] _0425_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0487_ counter2\[13\] counter2\[12\] counter2\[11\] counter2\[10\] _0317_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_0556_ _0377_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_26_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_5_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0949__55 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0851__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0608_ counter5\[1\] counter5\[0\] counter5\[2\] _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0539_ _0362_ _0363_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0803__176 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0946__58 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0874__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_0__f_clk clknet_0_clk clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0890_ net101 clknet_leaf_23_clk counter2\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0747__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0873_ net118 clknet_leaf_25_clk counter2\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_30_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0942_ net62 clknet_leaf_3_clk counter10\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_45_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0800__179 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0912__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0787_ net192 clknet_leaf_20_clk counter5\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0856_ net132 clknet_leaf_32_clk counter3\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0925_ net68 clknet_leaf_39_clk counter\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0935__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0710_ counter8\[1\] _0290_ counter8\[2\] _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0595__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0641_ counter10\[8\] _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__0808__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0572_ _0393_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0958__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_45_clk clknet_2_0__leaf_clk clknet_leaf_45_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0839_ _0002_ clknet_leaf_25_clk net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0908_ net85 clknet_leaf_42_clk counter\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_clk clknet_2_2__leaf_clk clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_27_clk clknet_2_3__leaf_clk clknet_leaf_27_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0624_ _0341_ _0425_ _0426_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0486_ counter2\[9\] counter2\[8\] counter2\[7\] counter2\[6\] _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_0555_ counter9\[26\] counter9\[25\] counter9\[23\] counter9\[24\] _0378_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__0780__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_18_clk clknet_2_1__leaf_clk clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_41_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0767__206 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_21_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1009__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0538_ counter7\[9\] counter7\[10\] counter7\[11\] counter7\[12\] _0363_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_7_clk clknet_2_1__leaf_clk clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0607_ _0409_ _0416_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0764__209 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0991__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0841__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0942__62 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_45_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0941_ net63 clknet_leaf_2_clk counter10\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0872_ net119 clknet_leaf_25_clk counter2\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0887__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0737__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0924_ net69 clknet_leaf_37_clk counter\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0786_ _0069_ clknet_leaf_27_clk counter5\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0855_ net133 clknet_leaf_43_clk counter3\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_44_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0640_ _0310_ _0314_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0571_ _0392_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0907_ net86 clknet_leaf_36_clk counter\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0838_ net146 clknet_leaf_7_clk counter4\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0769_ net204 clknet_leaf_45_clk counter6\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0902__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0554_ counter9\[22\] counter9\[21\] counter9\[20\] counter9\[19\] _0377_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_0623_ counter4\[0\] counter4\[1\] _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0485_ counter2\[5\] counter2\[4\] counter2\[3\] counter2\[2\] _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_38_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0948__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0537_ counter7\[13\] counter7\[14\] counter7\[15\] counter7\[16\] _0362_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0606_ counter6\[5\] _0414_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0773__200 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_14_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0631__A2 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0940_ net64 clknet_leaf_49_clk counter10\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0871_ net120 clknet_leaf_25_clk counter2\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0763__210 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_51_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0770__203 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0854_ net134 clknet_leaf_32_clk counter3\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0923_ net70 clknet_leaf_38_clk counter\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0785_ _0068_ clknet_leaf_30_clk counter5\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0831__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0589__A1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0760__213 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0570_ _0385_ _0387_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0837_ net147 clknet_leaf_7_clk counter4\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0906_ net87 clknet_leaf_38_clk counter\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0699_ _0376_ _0459_ _0461_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0768_ net205 clknet_leaf_46_clk counter6\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0727__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0877__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0967__47 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0622_ counter4\[0\] counter4\[1\] _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_0553_ counter9\[8\] _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0484_ _0310_ _0314_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0716__A1 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_43_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0536_ counter7\[25\] counter7\[24\] _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0605_ _0359_ _0414_ _0415_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0954__50 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0915__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0519_ counter5\[10\] counter5\[9\] counter5\[8\] counter5\[7\] _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_0951__53 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0938__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0870_ _0150_ clknet_leaf_25_clk counter2\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0999_ net24 clknet_leaf_16_clk counter8\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0760__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0853_ net135 clknet_leaf_43_clk counter3\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0922_ net71 clknet_leaf_37_clk counter\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0598__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0572__I _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0783__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0784_ _0067_ clknet_leaf_27_clk counter5\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_48_clk clknet_2_0__leaf_clk clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_39_clk clknet_2_2__leaf_clk clknet_leaf_39_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_clk_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0504__A2 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0836_ net148 clknet_leaf_8_clk counter4\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0905_ net88 clknet_leaf_40_clk counter\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0767_ net206 clknet_leaf_47_clk counter6\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0698_ _0472_ _0473_ _0474_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_2_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0621_ counter4\[0\] _0341_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0829__155 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0552_ counter8\[7\] _0375_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0821__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0483_ _0311_ _0312_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0836__148 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0819_ net165 clknet_leaf_5_clk counter4\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0844__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0994__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0604_ counter6\[4\] _0407_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0535_ counter7\[27\] counter7\[26\] counter7\[7\] counter7\[8\] _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0867__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0819__165 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_27_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0826__158 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_42_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0518_ counter5\[18\] counter5\[17\] counter5\[16\] counter5\[15\] _0345_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0607__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0998_ net25 clknet_leaf_18_clk counter8\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0909__84 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0905__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0816__168 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_27_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0921_ net72 clknet_leaf_38_clk counter\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0783_ _0066_ clknet_2_3__leaf_clk counter5\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0852_ net136 clknet_leaf_41_clk counter3\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0906__87 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0979__35 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0797__182 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0750__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0904_ net89 clknet_leaf_40_clk counter\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0835_ net149 clknet_leaf_7_clk counter4\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0697_ _0379_ _0383_ _0459_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0766_ net207 clknet_leaf_45_clk counter6\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0976__38 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_20_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0773__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0551_ _0370_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0620_ _0349_ _0419_ _0424_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0482_ counter\[12\] counter\[11\] counter\[9\] counter\[10\] _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_53_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0749_ net217 clknet_leaf_11_clk counter7\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0818_ net166 clknet_leaf_19_clk counter4\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0796__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0787__192 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0794__185 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_2_1__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0534_ counter6\[5\] _0359_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0603_ counter6\[4\] _0407_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_1_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0811__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0961__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0517_ counter5\[14\] counter5\[13\] counter5\[12\] counter5\[11\] _0344_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0834__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0791__188 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0832__152 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_13_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0857__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1008__15 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0997_ net26 clknet_leaf_18_clk counter8\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1012__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0747__219 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_41_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0920_ net73 clknet_leaf_38_clk counter\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1005__18 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0782_ _0065_ clknet_leaf_26_clk counter5\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0851_ net137 clknet_leaf_43_clk counter3\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0822__162 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0834_ net150 clknet_leaf_3_clk counter4\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0903_ net90 clknet_leaf_40_clk counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0696_ counter9\[6\] _0466_ _0458_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_0765_ net208 clknet_leaf_45_clk counter6\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0737__229 net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0902__91 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0723__B _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0918__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0550_ _0371_ _0372_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_7_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0481_ counter\[8\] counter\[7\] counter\[6\] counter\[5\] _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_19_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0817_ net167 clknet_leaf_5_clk counter4\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0748_ net218 clknet_leaf_10_clk counter7\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0679_ counter9\[1\] _0456_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_37_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0972__42 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0740__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0890__CLK clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0602_ _0359_ _0407_ _0413_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0533_ _0352_ _0355_ _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0763__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_clk clknet_2_1__leaf_clk clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0516_ counter5\[26\] counter5\[25\] counter5\[24\] counter5\[23\] _0343_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0543__A2 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_0_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0918__75 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0996_ net27 clknet_leaf_17_clk counter8\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0801__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0951__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0915__78 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0997__26 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_41_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0850_ net138 clknet_leaf_45_clk counter3\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0781_ _0004_ clknet_leaf_2_clk net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0824__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0974__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_1__f_clk clknet_0_clk clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0746__220 net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0979_ net35 clknet_leaf_30_clk counter9\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0994__29 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0847__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0997__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0833_ net151 clknet_leaf_3_clk counter4\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0902_ net91 clknet_leaf_36_clk counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1001__22 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1002__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0695_ counter9\[7\] _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0764_ net209 clknet_leaf_46_clk counter6\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_40_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0719__A2 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0480_ counter\[4\] counter\[3\] counter\[2\] counter\[27\] _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_66_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0736__230 net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0747_ net219 clknet_leaf_9_clk counter7\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0743__223 net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0816_ net168 clknet_leaf_18_clk counter4\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0678_ _0456_ _0461_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0750__216 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0859__129 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0601_ counter6\[2\] _0410_ counter6\[3\] _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0532_ _0356_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0908__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0561__A3 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0733__233 net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0515_ counter5\[22\] counter5\[21\] counter5\[20\] counter5\[19\] _0342_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_0740__226 net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0849__139 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0880__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0753__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0995_ net28 clknet_leaf_17_clk counter8\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0776__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0780_ net193 clknet_leaf_46_clk counter6\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0978_ net36 clknet_leaf_34_clk counter9\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0799__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0911__82 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0993__30 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0832_ net152 clknet_leaf_3_clk counter4\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0901_ net92 clknet_leaf_39_clk counter\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0763_ net210 clknet_leaf_46_clk counter6\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0694_ _0464_ _0471_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0941__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0814__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0964__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0746_ net220 clknet_leaf_9_clk counter7\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0815_ net169 clknet_leaf_6_clk counter4\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0981__33 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0677_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0837__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0987__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0531_ counter6\[9\] counter6\[8\] counter6\[7\] counter6\[6\] _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_11_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0600_ _0409_ _0412_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1014_ _0289_ clknet_leaf_13_clk counter7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0729_ _0014_ clknet_leaf_12_clk counter7\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0858__130 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_27_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0865__123 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0514_ counter4\[3\] _0341_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0994_ net29 clknet_leaf_17_clk counter8\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0848__140 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0924__69 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0855__133 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0862__126 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_18_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0870__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0977_ net37 clknet_leaf_30_clk counter9\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1010__13 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0743__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0893__CLK clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0900_ net93 clknet_leaf_39_clk counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0831_ net153 clknet_leaf_8_clk counter4\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0693_ counter9\[6\] _0470_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_0762_ net211 clknet_leaf_45_clk counter6\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0845__143 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0852__136 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0766__CLK clknet_leaf_45_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_50_clk clknet_2_0__leaf_clk clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0789__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0814_ _0096_ clknet_leaf_3_clk counter4\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_41_clk clknet_2_2__leaf_clk clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_14_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0745_ net221 clknet_leaf_10_clk counter7\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0676_ _0376_ _0459_ _0383_ _0379_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_32_clk clknet_2_2__leaf_clk clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_16_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0530_ counter6\[13\] counter6\[12\] counter6\[10\] counter6\[11\] _0356_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1013_ _0006_ clknet_leaf_48_clk net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_14_clk clknet_2_1__leaf_clk clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0728_ _0013_ clknet_leaf_11_clk counter7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0659_ counter10\[4\] _0447_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0954__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0513_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__0827__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0977__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0993_ net30 clknet_leaf_17_clk counter8\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1005__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0923__70 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_18_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0976_ net38 clknet_leaf_31_clk counter9\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0600__A1 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0920__73 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0830_ net154 clknet_leaf_4_clk counter4\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0692_ _0457_ _0458_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0761_ net212 clknet_leaf_4_clk counter6\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0959_ _0236_ clknet_leaf_36_clk counter9\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0860__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0813_ _0095_ clknet_leaf_2_clk counter4\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0744_ net222 clknet_leaf_8_clk counter7\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0675_ counter9\[7\] counter9\[6\] _0457_ _0458_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0733__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0513__I _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1012_ net11 clknet_leaf_14_clk counter8\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0756__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0727_ _0012_ clknet_leaf_13_clk counter7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0939__65 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0589_ _0367_ _0404_ _0405_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0658_ _0392_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0779__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0512_ _0333_ _0334_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0777__196 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0888__103 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0921__CLK clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0992_ _0268_ clknet_leaf_15_clk counter8\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0944__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0817__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0967__CLK clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0878__113 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0774__199 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0885__106 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0975_ net39 clknet_leaf_30_clk counter9\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0760_ net213 clknet_leaf_4_clk counter6\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0691_ _0466_ _0458_ _0464_ _0469_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0889_ net102 clknet_leaf_24_clk counter2\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0958_ _0235_ clknet_leaf_33_clk counter9\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0875__116 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_19_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0896__95 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_61_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0882__109 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0743_ net223 clknet_leaf_7_clk counter7\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0812_ _0094_ clknet_leaf_8_clk counter4\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0674_ counter9\[5\] counter9\[4\] _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0893__98 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1011_ net12 clknet_leaf_14_clk counter8\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0726_ _0011_ clknet_leaf_14_clk counter7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0588_ counter7\[5\] _0402_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0657_ _0392_ _0439_ _0446_ _0447_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_40_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0850__CLK clknet_leaf_45_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0872__119 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0511_ _0335_ _0336_ _0337_ _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0873__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0709_ counter8\[2\] counter8\[1\] _0290_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_38_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0896__CLK clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0746__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0991_ _0267_ clknet_leaf_15_clk counter8\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0769__CLK clknet_leaf_45_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0808__171 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0974_ net40 clknet_leaf_33_clk counter9\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0911__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0934__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0690_ counter9\[4\] _0466_ counter9\[5\] _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0780__193 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0891__100 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_52_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_44_clk clknet_2_0__leaf_clk clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0888_ net103 clknet_leaf_22_clk counter2\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0957_ _0234_ clknet_leaf_33_clk counter9\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0807__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0957__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_35_clk clknet_2_2__leaf_clk clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0805__174 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_26_clk clknet_2_3__leaf_clk clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0742_ net224 clknet_leaf_9_clk counter7\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0811_ _0093_ clknet_leaf_8_clk counter4\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0673_ counter9\[3\] counter9\[2\] counter9\[1\] counter9\[0\] _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_clk clknet_2_1__leaf_clk clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_19_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0881__110 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0948__56 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1010_ net13 clknet_leaf_13_clk counter8\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0725_ _0010_ clknet_leaf_14_clk counter7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1008__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_6_clk clknet_2_1__leaf_clk clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0656_ _0436_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0587_ counter7\[5\] _0402_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0802__177 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0945__59 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0510_ counter4\[7\] counter4\[6\] counter4\[5\] counter4\[4\] _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0630__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0639_ _0323_ _0434_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0708_ _0295_ _0296_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0871__120 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0990_ _0266_ clknet_leaf_17_clk counter8\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0840__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0990__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0973_ net41 clknet_leaf_32_clk counter9\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0736__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0886__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0769__204 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_52_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0899__94 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0759__CLK clknet_leaf_45_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0956_ _0233_ clknet_leaf_33_clk counter9\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0887_ net104 clknet_leaf_24_clk counter2\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0810_ _0003_ clknet_leaf_40_clk net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0741_ net225 clknet_leaf_9_clk counter7\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0672_ counter9\[0\] _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0939_ net65 clknet_leaf_1_clk counter10\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0924__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0759__214 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xclkbuf_2_2__f_clk clknet_0_clk clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0766__207 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0947__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0724_ counter7\[0\] _0398_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0586_ _0367_ _0402_ _0403_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0655_ counter10\[3\] _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_50_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0944__60 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_18_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0707_ counter8\[1\] _0290_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0638_ counter2\[1\] counter2\[0\] _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__0697__A2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0569_ _0388_ _0389_ _0390_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_57_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0941__63 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0792__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0972_ net42 clknet_leaf_32_clk counter9\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0830__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0955_ _0008_ clknet_leaf_15_clk net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0886_ net105 clknet_leaf_24_clk counter2\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0853__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0740_ net226 clknet_leaf_9_clk counter7\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0726__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0671_ _0385_ _0455_ _0443_ _0393_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__0876__CLK clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0869_ _0149_ clknet_leaf_25_clk counter2\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0938_ net66 clknet_leaf_1_clk counter10\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0749__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0899__CLK clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0723_ _0291_ _0293_ _0295_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0585_ counter7\[4\] _0395_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0654_ _0392_ _0443_ _0444_ _0445_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0772__201 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0914__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0706_ _0290_ _0295_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0637_ counter2\[0\] _0323_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0499_ counter3\[24\] counter3\[23\] counter3\[22\] counter3\[21\] _0328_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_0568_ counter10\[21\] counter10\[20\] counter10\[19\] counter10\[18\] _0390_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_53_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0937__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0762__211 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_17_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0971_ net43 clknet_leaf_32_clk counter9\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_47_clk clknet_2_0__leaf_clk clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0782__CLK clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_38_clk clknet_2_2__leaf_clk clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_clk clknet_2_3__leaf_clk clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0885_ net106 clknet_leaf_21_clk counter2\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0969__45 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0954_ net50 clknet_leaf_1_clk counter10\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0966__48 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0670_ _0435_ _0438_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_clk clknet_2_1__leaf_clk clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0799_ net180 clknet_leaf_18_clk counter5\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0868_ _0001_ clknet_leaf_38_clk net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0937_ net67 clknet_leaf_1_clk counter10\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0820__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0970__CLK clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0706__A2 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0722_ _0375_ _0304_ _0305_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_6_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0653_ counter10\[1\] _0441_ counter10\[2\] _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_8_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0584_ counter7\[4\] _0395_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0843__CLK clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0993__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0633__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0953__51 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_33_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0705_ _0294_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0636_ _0332_ _0433_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0950__54 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0567_ counter10\[17\] counter10\[16\] counter10\[15\] counter10\[14\] _0389_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_0498_ counter3\[25\] counter3\[26\] _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0739__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0889__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0619_ counter5\[4\] _0418_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0904__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0970_ net44 clknet_leaf_31_clk counter9\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0838__146 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0884_ net107 clknet_leaf_21_clk counter2\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0953_ net51 clknet_leaf_1_clk counter10\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_16_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_2_0__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0660__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0772__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0936_ _0214_ clknet_leaf_0_clk counter10\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0798_ net181 clknet_leaf_20_clk counter5\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0828__156 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0867_ net121 clknet_leaf_42_clk counter3\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0835__149 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0795__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0721_ counter8\[6\] _0302_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0583_ _0395_ _0397_ _0401_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0652_ counter10\[1\] _0441_ counter10\[2\] _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0919_ net74 clknet_leaf_38_clk counter\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0818__166 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0810__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0704_ _0291_ _0293_ _0374_ _0370_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_0825__159 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0960__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0635_ counter3\[2\] _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0566_ counter10\[13\] counter10\[12\] counter10\[11\] counter10\[10\] _0388_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_57_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0497_ counter3\[12\] counter3\[11\] counter3\[10\] counter3\[9\] _0326_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_53_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0833__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0983__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0618_ _0349_ _0418_ _0423_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0799__180 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0549_ counter8\[18\] counter8\[19\] counter8\[17\] counter8\[16\] _0373_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_0908__85 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1011__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0815__169 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_32_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0879__CLK clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0905__88 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_50_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0978__36 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0503__A4 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0952_ net52 clknet_leaf_2_clk counter10\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0883_ net108 clknet_leaf_21_clk counter2\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0789__190 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_9_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0796__183 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_28_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0975__39 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_23_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0917__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0866_ net122 clknet_leaf_44_clk counter3\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0935_ _0213_ clknet_leaf_1_clk counter10\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0797_ net182 clknet_leaf_18_clk counter5\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0720_ _0293_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0582_ counter7\[2\] _0394_ counter7\[3\] _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0651_ _0439_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_15_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0793__186 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0834__150 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_25_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0849_ net139 clknet_leaf_41_clk counter3\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0918_ net75 clknet_leaf_35_clk counter\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0762__CLK clknet_leaf_45_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0703_ counter8\[6\] counter8\[4\] counter8\[5\] _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_0749__217 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xclkbuf_leaf_10_clk clknet_2_1__leaf_clk clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0496_ counter3\[7\] counter3\[8\] counter3\[6\] counter3\[5\] _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_0634_ counter3\[1\] counter3\[0\] _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0565_ counter10\[27\] counter10\[26\] _0386_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0785__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0824__160 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_67_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0790__189 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0831__153 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_1007__16 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0617_ counter5\[3\] _0417_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0548_ counter8\[12\] counter8\[13\] counter8\[14\] counter8\[15\] _0372_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_0479_ _0306_ _0307_ _0308_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0739__227 net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0800__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0950__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1004__19 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0823__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_49_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0821__163 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0882_ net109 clknet_leaf_25_clk counter2\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0951_ net53 clknet_leaf_2_clk counter10\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0846__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0996__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0663__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0901__92 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1001__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0869__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0974__40 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0865_ net123 clknet_leaf_43_clk counter3\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0934_ _0212_ clknet_leaf_49_clk counter10\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0796_ net183 clknet_leaf_22_clk counter5\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0636__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0971__43 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_47_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0581_ _0398_ _0400_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0650_ _0393_ _0440_ _0442_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0848_ net140 clknet_leaf_43_clk counter3\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0779_ net194 clknet_leaf_48_clk counter6\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0917_ net76 clknet_leaf_35_clk counter\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0907__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0702_ counter8\[2\] counter8\[3\] counter8\[1\] counter8\[0\] _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_30_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0633_ _0332_ _0431_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0495_ counter3\[4\] counter3\[3\] counter3\[27\] _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0564_ counter10\[25\] counter10\[24\] counter10\[23\] counter10\[22\] _0386_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_14_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_29_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0917__76 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0999__24 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0616_ _0350_ _0417_ _0422_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0547_ counter8\[10\] counter8\[11\] counter8\[9\] counter8\[8\] _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_26_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0478_ counter\[26\] counter\[25\] counter\[1\] counter\[0\] _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__0752__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0914__79 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0996__27 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0775__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1003__20 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0745__221 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_41_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0798__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0881_ net110 clknet_leaf_26_clk counter2\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0950_ net54 clknet_leaf_2_clk counter10\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1000__23 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0940__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0813__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0795_ net184 clknet_leaf_22_clk counter5\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0963__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0864_ net124 clknet_leaf_44_clk counter3\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0933_ _0211_ clknet_leaf_49_clk counter10\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0735__231 net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0742__224 net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0836__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0986__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0580_ counter7\[2\] _0394_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0916_ net77 clknet_leaf_36_clk counter\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0778_ net195 clknet_leaf_48_clk counter6\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0847_ net141 clknet_leaf_33_clk counter3\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0859__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1014__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0701_ counter8\[7\] _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0632_ counter3\[1\] counter3\[0\] _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0563_ counter10\[9\] _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_0494_ counter2\[1\] _0323_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0732__234 net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_3__f_clk clknet_0_clk clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_58_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0546_ _0368_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0615_ counter5\[2\] _0420_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0477_ counter\[24\] counter\[23\] counter\[22\] counter\[21\] _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA_clkbuf_2_3__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0913__80 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_output8_I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0529_ _0353_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_13_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0910__83 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0880_ net111 clknet_leaf_24_clk counter2\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0742__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0892__CLK clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0983__31 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0765__CLK clknet_leaf_45_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0932_ _0210_ clknet_leaf_49_clk counter10\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_40_clk clknet_2_2__leaf_clk clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0867__121 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0794_ net185 clknet_leaf_22_clk counter5\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0863_ net125 clknet_leaf_44_clk counter3\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0980__34 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_28_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0788__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_31_clk clknet_2_3__leaf_clk clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_22_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_13_clk clknet_2_1__leaf_clk clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0915_ net78 clknet_leaf_36_clk counter\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0777_ net196 clknet_leaf_49_clk counter6\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0846_ net142 clknet_leaf_43_clk counter3\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0803__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0857__131 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0953__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0700_ counter8\[0\] _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0864__124 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0562_ _0384_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0631_ counter3\[0\] _0332_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_0493_ _0315_ _0316_ _0317_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0829_ net155 clknet_leaf_4_clk counter4\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0826__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0976__CLK clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0849__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0545_ counter8\[27\] counter8\[26\] counter8\[24\] counter8\[25\] _0369_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0614_ _0350_ _0420_ _0421_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0476_ counter\[16\] counter\[15\] counter\[13\] counter\[14\] _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1004__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0847__141 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0854__134 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1012__11 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0861__127 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0528_ counter6\[21\] counter6\[20\] counter6\[18\] counter6\[19\] _0354_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0648__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0844__144 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0851__137 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_12_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0862_ net126 clknet_leaf_44_clk counter3\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0931_ _0209_ clknet_leaf_50_clk counter10\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0793_ net186 clknet_leaf_16_clk counter5\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_27_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0732__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0882__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0845_ net143 clknet_leaf_43_clk counter3\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0914_ net79 clknet_leaf_37_clk counter\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0776_ net197 clknet_leaf_49_clk counter6\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0492_ _0318_ _0319_ _0320_ _0321_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_0561_ _0376_ _0379_ _0383_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_0630_ _0340_ _0429_ _0430_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0778__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0828_ net156 clknet_leaf_4_clk counter4\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0759_ net214 clknet_leaf_45_clk counter6\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0920__CLK clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0613_ counter5\[1\] counter5\[0\] _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0544_ counter8\[20\] counter8\[21\] counter8\[23\] counter8\[22\] _0368_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0475_ counter\[20\] counter\[19\] counter\[18\] counter\[17\] _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_53_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0943__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0922__71 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0816__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0966__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0527_ counter6\[17\] counter6\[16\] counter6\[14\] counter6\[15\] _0353_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0666__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0839__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput1 net1 cout1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0648__A2 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0792_ net187 clknet_leaf_30_clk counter5\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0861_ net127 clknet_leaf_5_clk counter3\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0930_ _0208_ clknet_leaf_50_clk counter10\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0779__194 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0775_ net198 clknet_leaf_49_clk counter6\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0844_ net144 clknet_leaf_42_clk counter3\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0913_ net80 clknet_leaf_36_clk counter\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0938__66 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_11_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_26_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0491_ counter2\[17\] counter2\[16\] counter2\[15\] counter2\[14\] _0321_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_0560_ _0380_ _0381_ _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0827_ net157 clknet_leaf_4_clk counter4\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0758_ _0042_ clknet_leaf_48_clk counter6\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0689_ _0461_ _0468_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0872__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0887__104 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0776__197 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0745__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0612_ counter5\[1\] counter5\[0\] _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0543_ counter7\[6\] _0367_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0895__CLK clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0768__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0877__114 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0526_ counter6\[27\] counter6\[26\] _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1009_ net14 clknet_leaf_14_clk counter8\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0884__107 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0910__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput2 net2 cout10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xclkbuf_leaf_43_clk clknet_2_2__leaf_clk clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0933__CLK clknet_leaf_49_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0509_ counter4\[11\] counter4\[10\] counter4\[9\] counter4\[8\] _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_34_clk clknet_2_2__leaf_clk clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0806__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0956__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0895__96 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xclkbuf_leaf_25_clk clknet_2_3__leaf_clk clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0791_ net188 clknet_leaf_19_clk counter5\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0860_ net128 clknet_leaf_19_clk counter3\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0874__117 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_51_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_16_clk clknet_2_1__leaf_clk clknet_leaf_16_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0989_ _0265_ clknet_leaf_16_clk counter8\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0829__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0979__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0892__99 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_42_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0912_ net81 clknet_leaf_36_clk counter\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0774_ net199 clknet_leaf_42_clk counter6\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0843_ net145 clknet_leaf_42_clk counter3\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0711__A2 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_5_clk clknet_2_0__leaf_clk clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1007__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0490_ counter2\[21\] counter2\[20\] counter2\[19\] counter2\[18\] _0320_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0705__I _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0826_ net158 clknet_leaf_6_clk counter4\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0688_ counter9\[4\] _0457_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_0757_ _0041_ clknet_leaf_48_clk counter6\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0542_ _0361_ _0364_ _0366_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0611_ counter5\[0\] _0350_ _0419_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_10_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0809_ net170 clknet_leaf_20_clk counter5\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_25_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0807__172 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0525_ counter6\[25\] counter6\[24\] counter6\[23\] counter6\[22\] _0351_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1008_ net15 clknet_leaf_14_clk counter8\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0735__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput3 net3 cout2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0508_ counter4\[18\] counter4\[19\] counter4\[17\] counter4\[16\] _0336_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0890__101 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0758__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0790_ net189 clknet_leaf_19_clk counter5\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0804__175 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0988_ _0264_ clknet_leaf_15_clk counter8\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0493__A2 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0947__57 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0923__CLK clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0842_ _0123_ clknet_leaf_40_clk counter3\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0911_ net82 clknet_leaf_36_clk counter\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0880__111 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0773_ net200 clknet_leaf_41_clk counter6\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0946__CLK clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0801__178 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0819__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0969__CLK clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0825_ net159 clknet_leaf_6_clk counter4\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0687_ _0466_ _0464_ _0467_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_0756_ _0040_ clknet_leaf_48_clk counter6\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0610_ counter5\[4\] _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_0541_ counter7\[21\] counter7\[22\] counter7\[23\] _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0791__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0808_ net171 clknet_leaf_30_clk counter5\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0739_ net227 clknet_leaf_10_clk counter7\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0524_ counter5\[4\] _0350_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1007_ net16 clknet_leaf_13_clk counter8\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput4 net4 cout3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_24_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0768__205 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_8_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0507_ counter4\[14\] counter4\[15\] counter4\[12\] counter4\[13\] _0335_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_27_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0852__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0987_ _0263_ clknet_leaf_22_clk counter8\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0725__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0875__CLK clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0772_ net201 clknet_leaf_41_clk counter6\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0841_ _0122_ clknet_leaf_40_clk counter3\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0765__208 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_0910_ net83 clknet_leaf_36_clk counter\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0748__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0898__CLK clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0943__61 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_21_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0824_ net160 clknet_leaf_6_clk counter4\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0755_ _0039_ clknet_leaf_47_clk counter6\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0686_ counter9\[3\] _0463_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0913__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0940__64 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_43_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0540_ counter7\[17\] counter7\[18\] counter7\[19\] counter7\[20\] _0365_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_3_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0738_ net228 clknet_leaf_7_clk counter7\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0807_ net172 clknet_leaf_30_clk counter5\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0669_ _0435_ _0438_ _0443_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0809__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0959__CLK clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0523_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1006_ net17 clknet_leaf_14_clk counter8\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_46_clk clknet_2_0__leaf_clk clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_41_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_37_clk clknet_2_2__leaf_clk clknet_leaf_37_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_53_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput5 net5 cout4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__0781__CLK clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0506_ counter4\[27\] counter4\[26\] counter4\[24\] counter4\[25\] _0334_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0986_ _0262_ clknet_leaf_15_clk counter8\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_8_clk clknet_2_1__leaf_clk clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_8_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0714__A2 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0650__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_23_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_38_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0771_ net202 clknet_leaf_47_clk counter6\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0840_ _0121_ clknet_leaf_42_clk counter3\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0969_ net45 clknet_leaf_31_clk counter9\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0992__CLK clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0842__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0771__202 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_9_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0823_ net161 clknet_leaf_6_clk counter4\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0685_ _0457_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0865__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0754_ _0038_ clknet_leaf_41_clk counter6\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0888__CLK clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0738__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0737_ net229 clknet_leaf_7_clk counter7\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0806_ net173 clknet_leaf_30_clk counter5\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0668_ _0448_ _0443_ _0454_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0599_ counter6\[2\] _0410_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0761__212 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0522_ _0342_ _0343_ _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0903__CLK clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1005_ net18 clknet_leaf_14_clk counter8\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput6 net6 cout5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_31_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0926__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0968__46 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0505_ counter4\[22\] counter4\[23\] counter4\[21\] counter4\[20\] _0333_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

