VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO divider
  CLASS BLOCK ;
  FOREIGN divider ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 218.400 4.000 218.960 ;
    END
  END clk
  PIN cout1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 26.880 299.000 27.440 ;
    END
  END cout1
  PIN cout10
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END cout10
  PIN cout2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.280 296.000 245.840 299.000 ;
    END
  END cout2
  PIN cout3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 1.000 218.960 4.000 ;
    END
  END cout3
  PIN cout4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 107.520 4.000 108.080 ;
    END
  END cout4
  PIN cout5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 245.280 299.000 245.840 ;
    END
  END cout5
  PIN cout6
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 1.000 108.080 4.000 ;
    END
  END cout6
  PIN cout7
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 296.000 27.440 299.000 ;
    END
  END cout7
  PIN cout8
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 296.000 134.960 299.000 ;
    END
  END cout8
  PIN cout9
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 134.400 299.000 134.960 ;
    END
  END cout9
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 283.210 ;
      LAYER Metal2 ;
        RECT 0.140 295.700 26.580 296.000 ;
        RECT 27.740 295.700 134.100 296.000 ;
        RECT 135.260 295.700 244.980 296.000 ;
        RECT 246.140 295.700 286.020 296.000 ;
        RECT 0.140 4.300 286.020 295.700 ;
        RECT 0.860 4.000 107.220 4.300 ;
        RECT 108.380 4.000 218.100 4.300 ;
        RECT 219.260 4.000 286.020 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 246.140 296.000 282.380 ;
        RECT 0.090 244.980 295.700 246.140 ;
        RECT 0.090 219.260 296.000 244.980 ;
        RECT 0.090 218.100 0.700 219.260 ;
        RECT 4.300 218.100 296.000 219.260 ;
        RECT 0.090 135.260 296.000 218.100 ;
        RECT 0.090 134.100 295.700 135.260 ;
        RECT 0.090 108.380 296.000 134.100 ;
        RECT 0.090 107.220 0.700 108.380 ;
        RECT 4.300 107.220 296.000 108.380 ;
        RECT 0.090 27.740 296.000 107.220 ;
        RECT 0.090 26.580 295.700 27.740 ;
        RECT 0.090 15.540 296.000 26.580 ;
  END
END divider
END LIBRARY

