magic
tech gf180mcuC
magscale 1 5
timestamp 1670270216
<< obsm1 >>
rect 672 1538 29288 28321
<< metal2 >>
rect 2688 29600 2744 29900
rect 13440 29600 13496 29900
rect 24528 29600 24584 29900
rect 0 100 56 400
rect 10752 100 10808 400
rect 21840 100 21896 400
<< obsm2 >>
rect 14 29570 2658 29600
rect 2774 29570 13410 29600
rect 13526 29570 24498 29600
rect 24614 29570 28602 29600
rect 14 430 28602 29570
rect 86 400 10722 430
rect 10838 400 21810 430
rect 21926 400 28602 430
<< metal3 >>
rect 29600 24528 29900 24584
rect 100 21840 400 21896
rect 29600 13440 29900 13496
rect 100 10752 400 10808
rect 29600 2688 29900 2744
<< obsm3 >>
rect 9 24614 29600 28238
rect 9 24498 29570 24614
rect 9 21926 29600 24498
rect 9 21810 70 21926
rect 430 21810 29600 21926
rect 9 13526 29600 21810
rect 9 13410 29570 13526
rect 9 10838 29600 13410
rect 9 10722 70 10838
rect 430 10722 29600 10838
rect 9 2774 29600 10722
rect 9 2658 29570 2774
rect 9 1554 29600 2658
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
rect 25264 1538 25424 28254
<< labels >>
rlabel metal3 s 100 21840 400 21896 6 clk
port 1 nsew signal input
rlabel metal3 s 29600 2688 29900 2744 6 cout1
port 2 nsew signal output
rlabel metal2 s 0 100 56 400 6 cout10
port 3 nsew signal output
rlabel metal2 s 24528 29600 24584 29900 6 cout2
port 4 nsew signal output
rlabel metal2 s 21840 100 21896 400 6 cout3
port 5 nsew signal output
rlabel metal3 s 100 10752 400 10808 6 cout4
port 6 nsew signal output
rlabel metal3 s 29600 24528 29900 24584 6 cout5
port 7 nsew signal output
rlabel metal2 s 10752 100 10808 400 6 cout6
port 8 nsew signal output
rlabel metal2 s 2688 29600 2744 29900 6 cout7
port 9 nsew signal output
rlabel metal2 s 13440 29600 13496 29900 6 cout8
port 10 nsew signal output
rlabel metal3 s 29600 13440 29900 13496 6 cout9
port 11 nsew signal output
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 12 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 12 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 13 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 28254 6 vss
port 13 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1442356
string GDS_FILE /home/urielcho/Proyectos_caravel/gf180nm/divider/openlane/divider/runs/22_12_05_13_55/results/signoff/divider.magic.gds
string GDS_START 156512
<< end >>

