magic
tech gf180mcuC
magscale 1 10
timestamp 1670270215
<< metal1 >>
rect 5394 56590 5406 56642
rect 5458 56639 5470 56642
rect 6402 56639 6414 56642
rect 5458 56593 6414 56639
rect 5458 56590 5470 56593
rect 6402 56590 6414 56593
rect 6466 56590 6478 56642
rect 26898 56590 26910 56642
rect 26962 56639 26974 56642
rect 27794 56639 27806 56642
rect 26962 56593 27806 56639
rect 26962 56590 26974 56593
rect 27794 56590 27806 56593
rect 27858 56590 27870 56642
rect 49074 56590 49086 56642
rect 49138 56639 49150 56642
rect 49970 56639 49982 56642
rect 49138 56593 49982 56639
rect 49138 56590 49150 56593
rect 49970 56590 49982 56593
rect 50034 56590 50046 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 5070 56082 5122 56094
rect 5730 56030 5742 56082
rect 5794 56030 5806 56082
rect 27234 56030 27246 56082
rect 27298 56030 27310 56082
rect 49298 56030 49310 56082
rect 49362 56030 49374 56082
rect 5070 56018 5122 56030
rect 6402 55918 6414 55970
rect 6466 55918 6478 55970
rect 27794 55918 27806 55970
rect 27858 55918 27870 55970
rect 49970 55918 49982 55970
rect 50034 55918 50046 55970
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 8318 52162 8370 52174
rect 8318 52098 8370 52110
rect 9102 52162 9154 52174
rect 9102 52098 9154 52110
rect 8430 51938 8482 51950
rect 8430 51874 8482 51886
rect 8542 51938 8594 51950
rect 8542 51874 8594 51886
rect 19518 51938 19570 51950
rect 19518 51874 19570 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 41582 51490 41634 51502
rect 19282 51438 19294 51490
rect 19346 51438 19358 51490
rect 41582 51426 41634 51438
rect 9774 51378 9826 51390
rect 8978 51326 8990 51378
rect 9042 51326 9054 51378
rect 18498 51326 18510 51378
rect 18562 51326 18574 51378
rect 33954 51326 33966 51378
rect 34018 51326 34030 51378
rect 45938 51326 45950 51378
rect 46002 51326 46014 51378
rect 49522 51326 49534 51378
rect 49586 51326 49598 51378
rect 9774 51314 9826 51326
rect 13246 51266 13298 51278
rect 21982 51266 22034 51278
rect 4946 51214 4958 51266
rect 5010 51214 5022 51266
rect 21410 51214 21422 51266
rect 21474 51214 21486 51266
rect 13246 51202 13298 51214
rect 21982 51202 22034 51214
rect 26238 51266 26290 51278
rect 37438 51266 37490 51278
rect 53006 51266 53058 51278
rect 34738 51214 34750 51266
rect 34802 51214 34814 51266
rect 36866 51214 36878 51266
rect 36930 51214 36942 51266
rect 46610 51214 46622 51266
rect 46674 51214 46686 51266
rect 48738 51214 48750 51266
rect 48802 51214 48814 51266
rect 50306 51214 50318 51266
rect 50370 51214 50382 51266
rect 52434 51214 52446 51266
rect 52498 51214 52510 51266
rect 26238 51202 26290 51214
rect 37438 51202 37490 51214
rect 53006 51202 53058 51214
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 2034 50654 2046 50706
rect 2098 50654 2110 50706
rect 4162 50654 4174 50706
rect 4226 50654 4238 50706
rect 9426 50654 9438 50706
rect 9490 50654 9502 50706
rect 12898 50654 12910 50706
rect 12962 50654 12974 50706
rect 13682 50654 13694 50706
rect 13746 50654 13758 50706
rect 27234 50654 27246 50706
rect 27298 50654 27310 50706
rect 40786 50654 40798 50706
rect 40850 50654 40862 50706
rect 42914 50654 42926 50706
rect 42978 50654 42990 50706
rect 4946 50542 4958 50594
rect 5010 50542 5022 50594
rect 6514 50542 6526 50594
rect 6578 50542 6590 50594
rect 10098 50542 10110 50594
rect 10162 50542 10174 50594
rect 16594 50542 16606 50594
rect 16658 50542 16670 50594
rect 24434 50542 24446 50594
rect 24498 50542 24510 50594
rect 40002 50542 40014 50594
rect 40066 50542 40078 50594
rect 17054 50482 17106 50494
rect 34862 50482 34914 50494
rect 7298 50430 7310 50482
rect 7362 50430 7374 50482
rect 10770 50430 10782 50482
rect 10834 50430 10846 50482
rect 15810 50430 15822 50482
rect 15874 50430 15886 50482
rect 25106 50430 25118 50482
rect 25170 50430 25182 50482
rect 17054 50418 17106 50430
rect 34862 50418 34914 50430
rect 39454 50482 39506 50494
rect 39454 50418 39506 50430
rect 50318 50482 50370 50494
rect 50318 50418 50370 50430
rect 54238 50482 54290 50494
rect 54238 50418 54290 50430
rect 21646 50370 21698 50382
rect 21646 50306 21698 50318
rect 27694 50370 27746 50382
rect 27694 50306 27746 50318
rect 37662 50370 37714 50382
rect 37662 50306 37714 50318
rect 48974 50370 49026 50382
rect 48974 50306 49026 50318
rect 53342 50370 53394 50382
rect 53342 50306 53394 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 8654 50034 8706 50046
rect 8654 49970 8706 49982
rect 9886 50034 9938 50046
rect 9886 49970 9938 49982
rect 11678 50034 11730 50046
rect 11678 49970 11730 49982
rect 23326 50034 23378 50046
rect 23326 49970 23378 49982
rect 42702 50034 42754 50046
rect 42702 49970 42754 49982
rect 47630 50034 47682 50046
rect 47630 49970 47682 49982
rect 9774 49922 9826 49934
rect 9774 49858 9826 49870
rect 12462 49922 12514 49934
rect 12462 49858 12514 49870
rect 12686 49922 12738 49934
rect 12686 49858 12738 49870
rect 13918 49922 13970 49934
rect 13918 49858 13970 49870
rect 16382 49922 16434 49934
rect 25790 49922 25842 49934
rect 20738 49870 20750 49922
rect 20802 49870 20814 49922
rect 16382 49858 16434 49870
rect 25790 49858 25842 49870
rect 41694 49922 41746 49934
rect 41694 49858 41746 49870
rect 47742 49922 47794 49934
rect 47742 49858 47794 49870
rect 8318 49810 8370 49822
rect 4274 49758 4286 49810
rect 4338 49758 4350 49810
rect 8318 49746 8370 49758
rect 8654 49810 8706 49822
rect 8654 49746 8706 49758
rect 8990 49810 9042 49822
rect 42254 49810 42306 49822
rect 43486 49810 43538 49822
rect 10098 49758 10110 49810
rect 10162 49758 10174 49810
rect 11890 49758 11902 49810
rect 11954 49758 11966 49810
rect 13346 49758 13358 49810
rect 13410 49758 13422 49810
rect 19954 49758 19966 49810
rect 20018 49758 20030 49810
rect 27682 49758 27694 49810
rect 27746 49758 27758 49810
rect 36866 49758 36878 49810
rect 36930 49758 36942 49810
rect 42802 49758 42814 49810
rect 42866 49758 42878 49810
rect 43250 49758 43262 49810
rect 43314 49758 43326 49810
rect 46946 49758 46958 49810
rect 47010 49758 47022 49810
rect 51090 49758 51102 49810
rect 51154 49758 51166 49810
rect 56130 49758 56142 49810
rect 56194 49758 56206 49810
rect 8990 49746 9042 49758
rect 42254 49746 42306 49758
rect 43486 49746 43538 49758
rect 24894 49698 24946 49710
rect 26462 49698 26514 49710
rect 4946 49646 4958 49698
rect 5010 49646 5022 49698
rect 7074 49646 7086 49698
rect 7138 49646 7150 49698
rect 12786 49646 12798 49698
rect 12850 49646 12862 49698
rect 22866 49646 22878 49698
rect 22930 49646 22942 49698
rect 25666 49646 25678 49698
rect 25730 49646 25742 49698
rect 24894 49634 24946 49646
rect 26462 49634 26514 49646
rect 27134 49698 27186 49710
rect 30942 49698 30994 49710
rect 28354 49646 28366 49698
rect 28418 49646 28430 49698
rect 30482 49646 30494 49698
rect 30546 49646 30558 49698
rect 37874 49646 37886 49698
rect 37938 49646 37950 49698
rect 44034 49646 44046 49698
rect 44098 49646 44110 49698
rect 46162 49646 46174 49698
rect 46226 49646 46238 49698
rect 51874 49646 51886 49698
rect 51938 49646 51950 49698
rect 54002 49646 54014 49698
rect 54066 49646 54078 49698
rect 55346 49646 55358 49698
rect 55410 49646 55422 49698
rect 27134 49634 27186 49646
rect 30942 49634 30994 49646
rect 11566 49586 11618 49598
rect 11566 49522 11618 49534
rect 13582 49586 13634 49598
rect 13582 49522 13634 49534
rect 13806 49586 13858 49598
rect 13806 49522 13858 49534
rect 24782 49586 24834 49598
rect 24782 49522 24834 49534
rect 26014 49586 26066 49598
rect 47518 49586 47570 49598
rect 42914 49534 42926 49586
rect 42978 49534 42990 49586
rect 26014 49522 26066 49534
rect 47518 49522 47570 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 12574 49250 12626 49262
rect 12574 49186 12626 49198
rect 22094 49250 22146 49262
rect 22094 49186 22146 49198
rect 22318 49250 22370 49262
rect 22318 49186 22370 49198
rect 28366 49250 28418 49262
rect 28366 49186 28418 49198
rect 45838 49250 45890 49262
rect 45838 49186 45890 49198
rect 21870 49138 21922 49150
rect 36318 49138 36370 49150
rect 15138 49086 15150 49138
rect 15202 49086 15214 49138
rect 17266 49086 17278 49138
rect 17330 49086 17342 49138
rect 20738 49086 20750 49138
rect 20802 49086 20814 49138
rect 22978 49086 22990 49138
rect 23042 49086 23054 49138
rect 21870 49074 21922 49086
rect 36318 49074 36370 49086
rect 36766 49138 36818 49150
rect 37538 49086 37550 49138
rect 37602 49086 37614 49138
rect 39666 49086 39678 49138
rect 39730 49086 39742 49138
rect 41794 49086 41806 49138
rect 41858 49086 41870 49138
rect 43922 49086 43934 49138
rect 43986 49086 43998 49138
rect 52434 49086 52446 49138
rect 52498 49086 52510 49138
rect 56466 49086 56478 49138
rect 56530 49086 56542 49138
rect 36766 49074 36818 49086
rect 7310 49026 7362 49038
rect 7310 48962 7362 48974
rect 7534 49026 7586 49038
rect 7534 48962 7586 48974
rect 12350 49026 12402 49038
rect 26350 49026 26402 49038
rect 14354 48974 14366 49026
rect 14418 48974 14430 49026
rect 17938 48974 17950 49026
rect 18002 48974 18014 49026
rect 21634 48974 21646 49026
rect 21698 48974 21710 49026
rect 25890 48974 25902 49026
rect 25954 48974 25966 49026
rect 12350 48962 12402 48974
rect 26350 48962 26402 48974
rect 26686 49026 26738 49038
rect 26686 48962 26738 48974
rect 30270 49026 30322 49038
rect 30930 48974 30942 49026
rect 30994 48974 31006 49026
rect 40338 48974 40350 49026
rect 40402 48974 40414 49026
rect 41010 48974 41022 49026
rect 41074 48974 41086 49026
rect 45826 48974 45838 49026
rect 45890 48974 45902 49026
rect 49522 48974 49534 49026
rect 49586 48974 49598 49026
rect 53554 48974 53566 49026
rect 53618 48974 53630 49026
rect 30270 48962 30322 48974
rect 8766 48914 8818 48926
rect 26574 48914 26626 48926
rect 18610 48862 18622 48914
rect 18674 48862 18686 48914
rect 25106 48862 25118 48914
rect 25170 48862 25182 48914
rect 8766 48850 8818 48862
rect 26574 48850 26626 48862
rect 27022 48914 27074 48926
rect 27022 48850 27074 48862
rect 28702 48914 28754 48926
rect 28702 48850 28754 48862
rect 30046 48914 30098 48926
rect 30046 48850 30098 48862
rect 45502 48914 45554 48926
rect 45502 48850 45554 48862
rect 48974 48914 49026 48926
rect 56926 48914 56978 48926
rect 50306 48862 50318 48914
rect 50370 48862 50382 48914
rect 54338 48862 54350 48914
rect 54402 48862 54414 48914
rect 48974 48850 49026 48862
rect 56926 48850 56978 48862
rect 8542 48802 8594 48814
rect 7858 48750 7870 48802
rect 7922 48750 7934 48802
rect 8542 48738 8594 48750
rect 8654 48802 8706 48814
rect 22206 48802 22258 48814
rect 12898 48750 12910 48802
rect 12962 48750 12974 48802
rect 8654 48738 8706 48750
rect 22206 48738 22258 48750
rect 27806 48802 27858 48814
rect 27806 48738 27858 48750
rect 28478 48802 28530 48814
rect 28478 48738 28530 48750
rect 33854 48802 33906 48814
rect 33854 48738 33906 48750
rect 35198 48802 35250 48814
rect 35198 48738 35250 48750
rect 47182 48802 47234 48814
rect 47182 48738 47234 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 18734 48466 18786 48478
rect 18734 48402 18786 48414
rect 20974 48466 21026 48478
rect 20974 48402 21026 48414
rect 24670 48466 24722 48478
rect 24670 48402 24722 48414
rect 36990 48466 37042 48478
rect 36990 48402 37042 48414
rect 41470 48466 41522 48478
rect 41470 48402 41522 48414
rect 7310 48354 7362 48366
rect 7310 48290 7362 48302
rect 8542 48354 8594 48366
rect 8542 48290 8594 48302
rect 24446 48354 24498 48366
rect 24446 48290 24498 48302
rect 32510 48354 32562 48366
rect 44718 48354 44770 48366
rect 34402 48302 34414 48354
rect 34466 48302 34478 48354
rect 32510 48290 32562 48302
rect 44718 48290 44770 48302
rect 48078 48354 48130 48366
rect 48078 48290 48130 48302
rect 7422 48242 7474 48254
rect 7422 48178 7474 48190
rect 7646 48242 7698 48254
rect 7646 48178 7698 48190
rect 9662 48242 9714 48254
rect 9662 48178 9714 48190
rect 12574 48242 12626 48254
rect 12574 48178 12626 48190
rect 12798 48242 12850 48254
rect 12798 48178 12850 48190
rect 13134 48242 13186 48254
rect 24334 48242 24386 48254
rect 48750 48242 48802 48254
rect 13906 48190 13918 48242
rect 13970 48190 13982 48242
rect 27346 48190 27358 48242
rect 27410 48190 27422 48242
rect 32722 48190 32734 48242
rect 32786 48190 32798 48242
rect 33730 48190 33742 48242
rect 33794 48190 33806 48242
rect 37874 48190 37886 48242
rect 37938 48190 37950 48242
rect 44034 48190 44046 48242
rect 44098 48190 44110 48242
rect 49522 48190 49534 48242
rect 49586 48190 49598 48242
rect 13134 48178 13186 48190
rect 24334 48178 24386 48190
rect 48750 48178 48802 48190
rect 12910 48130 12962 48142
rect 17614 48130 17666 48142
rect 8530 48078 8542 48130
rect 8594 48078 8606 48130
rect 14018 48078 14030 48130
rect 14082 48078 14094 48130
rect 12910 48066 12962 48078
rect 17614 48066 17666 48078
rect 25678 48130 25730 48142
rect 31714 48078 31726 48130
rect 31778 48078 31790 48130
rect 36530 48078 36542 48130
rect 36594 48078 36606 48130
rect 38658 48078 38670 48130
rect 38722 48078 38734 48130
rect 40786 48078 40798 48130
rect 40850 48078 40862 48130
rect 44482 48078 44494 48130
rect 44546 48078 44558 48130
rect 51538 48078 51550 48130
rect 51602 48078 51614 48130
rect 25678 48066 25730 48078
rect 7758 48018 7810 48030
rect 7758 47954 7810 47966
rect 8766 48018 8818 48030
rect 25790 48018 25842 48030
rect 14242 47966 14254 48018
rect 14306 47966 14318 48018
rect 8766 47954 8818 47966
rect 25790 47954 25842 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 37774 47682 37826 47694
rect 21634 47630 21646 47682
rect 21698 47630 21710 47682
rect 37774 47618 37826 47630
rect 38222 47682 38274 47694
rect 38222 47618 38274 47630
rect 7870 47570 7922 47582
rect 7870 47506 7922 47518
rect 22206 47570 22258 47582
rect 37998 47570 38050 47582
rect 24322 47518 24334 47570
rect 24386 47518 24398 47570
rect 27906 47518 27918 47570
rect 27970 47518 27982 47570
rect 28802 47518 28814 47570
rect 28866 47518 28878 47570
rect 34626 47518 34638 47570
rect 34690 47518 34702 47570
rect 36754 47518 36766 47570
rect 36818 47518 36830 47570
rect 45490 47518 45502 47570
rect 45554 47518 45566 47570
rect 47954 47518 47966 47570
rect 48018 47518 48030 47570
rect 50082 47518 50094 47570
rect 50146 47518 50158 47570
rect 22206 47506 22258 47518
rect 37998 47506 38050 47518
rect 7646 47458 7698 47470
rect 7646 47394 7698 47406
rect 8654 47458 8706 47470
rect 8654 47394 8706 47406
rect 8878 47458 8930 47470
rect 8878 47394 8930 47406
rect 9102 47458 9154 47470
rect 12686 47458 12738 47470
rect 12226 47406 12238 47458
rect 12290 47406 12302 47458
rect 9102 47394 9154 47406
rect 12686 47394 12738 47406
rect 12798 47458 12850 47470
rect 21982 47458 22034 47470
rect 30718 47458 30770 47470
rect 31614 47458 31666 47470
rect 14130 47406 14142 47458
rect 14194 47406 14206 47458
rect 23202 47406 23214 47458
rect 23266 47406 23278 47458
rect 24210 47406 24222 47458
rect 24274 47406 24286 47458
rect 25106 47406 25118 47458
rect 25170 47406 25182 47458
rect 31042 47406 31054 47458
rect 31106 47406 31118 47458
rect 12798 47394 12850 47406
rect 21982 47394 22034 47406
rect 30718 47394 30770 47406
rect 31614 47394 31666 47406
rect 32174 47458 32226 47470
rect 33842 47406 33854 47458
rect 33906 47406 33918 47458
rect 37538 47406 37550 47458
rect 37602 47406 37614 47458
rect 47170 47406 47182 47458
rect 47234 47406 47246 47458
rect 54002 47406 54014 47458
rect 54066 47406 54078 47458
rect 55122 47406 55134 47458
rect 55186 47406 55198 47458
rect 32174 47394 32226 47406
rect 8430 47346 8482 47358
rect 8430 47282 8482 47294
rect 10110 47346 10162 47358
rect 10110 47282 10162 47294
rect 10446 47346 10498 47358
rect 23438 47346 23490 47358
rect 28478 47346 28530 47358
rect 12450 47294 12462 47346
rect 12514 47294 12526 47346
rect 16818 47294 16830 47346
rect 16882 47294 16894 47346
rect 24098 47294 24110 47346
rect 24162 47294 24174 47346
rect 25778 47294 25790 47346
rect 25842 47294 25854 47346
rect 10446 47282 10498 47294
rect 23438 47282 23490 47294
rect 28478 47282 28530 47294
rect 28702 47346 28754 47358
rect 28702 47282 28754 47294
rect 29486 47346 29538 47358
rect 29486 47282 29538 47294
rect 30830 47346 30882 47358
rect 30830 47282 30882 47294
rect 31838 47346 31890 47358
rect 31838 47282 31890 47294
rect 38334 47346 38386 47358
rect 38334 47282 38386 47294
rect 39118 47346 39170 47358
rect 39118 47282 39170 47294
rect 45614 47346 45666 47358
rect 45614 47282 45666 47294
rect 45838 47346 45890 47358
rect 45838 47282 45890 47294
rect 52110 47346 52162 47358
rect 53442 47294 53454 47346
rect 53506 47294 53518 47346
rect 55010 47294 55022 47346
rect 55074 47294 55086 47346
rect 52110 47282 52162 47294
rect 9214 47234 9266 47246
rect 7298 47182 7310 47234
rect 7362 47182 7374 47234
rect 9214 47170 9266 47182
rect 11902 47234 11954 47246
rect 11902 47170 11954 47182
rect 19518 47234 19570 47246
rect 19518 47170 19570 47182
rect 20750 47234 20802 47246
rect 31950 47234 32002 47246
rect 30258 47182 30270 47234
rect 30322 47182 30334 47234
rect 20750 47170 20802 47182
rect 31950 47170 32002 47182
rect 50542 47234 50594 47246
rect 50542 47170 50594 47182
rect 52670 47234 52722 47246
rect 54002 47182 54014 47234
rect 54066 47182 54078 47234
rect 52670 47170 52722 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 17614 46898 17666 46910
rect 17614 46834 17666 46846
rect 37102 46898 37154 46910
rect 37102 46834 37154 46846
rect 47182 46898 47234 46910
rect 47182 46834 47234 46846
rect 54574 46898 54626 46910
rect 54574 46834 54626 46846
rect 3502 46786 3554 46798
rect 8990 46786 9042 46798
rect 5730 46734 5742 46786
rect 5794 46734 5806 46786
rect 3502 46722 3554 46734
rect 8990 46722 9042 46734
rect 16942 46786 16994 46798
rect 16942 46722 16994 46734
rect 24670 46786 24722 46798
rect 24670 46722 24722 46734
rect 25678 46786 25730 46798
rect 25678 46722 25730 46734
rect 27806 46786 27858 46798
rect 38334 46786 38386 46798
rect 29138 46734 29150 46786
rect 29202 46734 29214 46786
rect 41682 46734 41694 46786
rect 41746 46734 41758 46786
rect 42018 46734 42030 46786
rect 42082 46734 42094 46786
rect 45154 46734 45166 46786
rect 45218 46734 45230 46786
rect 48514 46734 48526 46786
rect 48578 46734 48590 46786
rect 27806 46722 27858 46734
rect 38334 46722 38386 46734
rect 8542 46674 8594 46686
rect 5058 46622 5070 46674
rect 5122 46622 5134 46674
rect 8542 46610 8594 46622
rect 8654 46674 8706 46686
rect 8654 46610 8706 46622
rect 8878 46674 8930 46686
rect 26014 46674 26066 46686
rect 9874 46622 9886 46674
rect 9938 46622 9950 46674
rect 16146 46622 16158 46674
rect 16210 46622 16222 46674
rect 18386 46622 18398 46674
rect 18450 46622 18462 46674
rect 8878 46610 8930 46622
rect 26014 46610 26066 46622
rect 27470 46674 27522 46686
rect 41582 46674 41634 46686
rect 28466 46622 28478 46674
rect 28530 46622 28542 46674
rect 27470 46610 27522 46622
rect 41582 46610 41634 46622
rect 42366 46674 42418 46686
rect 46398 46674 46450 46686
rect 45826 46622 45838 46674
rect 45890 46622 45902 46674
rect 42366 46610 42418 46622
rect 46398 46610 46450 46622
rect 47070 46674 47122 46686
rect 47730 46622 47742 46674
rect 47794 46622 47806 46674
rect 48402 46622 48414 46674
rect 48466 46622 48478 46674
rect 51202 46622 51214 46674
rect 51266 46622 51278 46674
rect 47070 46610 47122 46622
rect 24782 46562 24834 46574
rect 7858 46510 7870 46562
rect 7922 46510 7934 46562
rect 10546 46510 10558 46562
rect 10610 46510 10622 46562
rect 12674 46510 12686 46562
rect 12738 46510 12750 46562
rect 13234 46510 13246 46562
rect 13298 46510 13310 46562
rect 15362 46510 15374 46562
rect 15426 46510 15438 46562
rect 22866 46510 22878 46562
rect 22930 46510 22942 46562
rect 24782 46498 24834 46510
rect 25790 46562 25842 46574
rect 25790 46498 25842 46510
rect 26126 46562 26178 46574
rect 26126 46498 26178 46510
rect 26910 46562 26962 46574
rect 31726 46562 31778 46574
rect 31266 46510 31278 46562
rect 31330 46510 31342 46562
rect 26910 46498 26962 46510
rect 31726 46498 31778 46510
rect 40798 46562 40850 46574
rect 49534 46562 49586 46574
rect 43026 46510 43038 46562
rect 43090 46510 43102 46562
rect 51986 46510 51998 46562
rect 52050 46510 52062 46562
rect 54114 46510 54126 46562
rect 54178 46510 54190 46562
rect 40798 46498 40850 46510
rect 49534 46498 49586 46510
rect 24894 46450 24946 46462
rect 24894 46386 24946 46398
rect 42590 46450 42642 46462
rect 42590 46386 42642 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 10334 46114 10386 46126
rect 10334 46050 10386 46062
rect 10782 46114 10834 46126
rect 10782 46050 10834 46062
rect 21758 46114 21810 46126
rect 29822 46114 29874 46126
rect 25890 46062 25902 46114
rect 25954 46062 25966 46114
rect 21758 46050 21810 46062
rect 29822 46050 29874 46062
rect 30158 46114 30210 46126
rect 30158 46050 30210 46062
rect 9214 46002 9266 46014
rect 2818 45950 2830 46002
rect 2882 45950 2894 46002
rect 4946 45950 4958 46002
rect 5010 45950 5022 46002
rect 9214 45938 9266 45950
rect 12910 46002 12962 46014
rect 12910 45938 12962 45950
rect 13582 46002 13634 46014
rect 21870 46002 21922 46014
rect 17378 45950 17390 46002
rect 17442 45950 17454 46002
rect 18722 45950 18734 46002
rect 18786 45950 18798 46002
rect 20850 45950 20862 46002
rect 20914 45950 20926 46002
rect 13582 45938 13634 45950
rect 21870 45938 21922 45950
rect 22878 46002 22930 46014
rect 48974 46002 49026 46014
rect 30818 45950 30830 46002
rect 30882 45950 30894 46002
rect 38322 45950 38334 46002
rect 38386 45950 38398 46002
rect 40450 45950 40462 46002
rect 40514 45950 40526 46002
rect 43922 45950 43934 46002
rect 43986 45950 43998 46002
rect 48402 45950 48414 46002
rect 48466 45950 48478 46002
rect 22878 45938 22930 45950
rect 48974 45938 49026 45950
rect 10446 45890 10498 45902
rect 2034 45838 2046 45890
rect 2098 45838 2110 45890
rect 10446 45826 10498 45838
rect 10670 45890 10722 45902
rect 22094 45890 22146 45902
rect 14466 45838 14478 45890
rect 14530 45838 14542 45890
rect 18050 45838 18062 45890
rect 18114 45838 18126 45890
rect 10670 45826 10722 45838
rect 22094 45826 22146 45838
rect 22318 45890 22370 45902
rect 22318 45826 22370 45838
rect 25566 45890 25618 45902
rect 29934 45890 29986 45902
rect 26114 45838 26126 45890
rect 26178 45838 26190 45890
rect 26786 45838 26798 45890
rect 26850 45838 26862 45890
rect 33618 45838 33630 45890
rect 33682 45838 33694 45890
rect 37650 45838 37662 45890
rect 37714 45838 37726 45890
rect 41010 45838 41022 45890
rect 41074 45838 41086 45890
rect 45602 45838 45614 45890
rect 45666 45838 45678 45890
rect 25566 45826 25618 45838
rect 29934 45826 29986 45838
rect 52110 45778 52162 45790
rect 15250 45726 15262 45778
rect 15314 45726 15326 45778
rect 25778 45726 25790 45778
rect 25842 45726 25854 45778
rect 32946 45726 32958 45778
rect 33010 45726 33022 45778
rect 41794 45726 41806 45778
rect 41858 45726 41870 45778
rect 46274 45726 46286 45778
rect 46338 45726 46350 45778
rect 52110 45714 52162 45726
rect 5630 45666 5682 45678
rect 5630 45602 5682 45614
rect 8094 45666 8146 45678
rect 8094 45602 8146 45614
rect 22206 45666 22258 45678
rect 22206 45602 22258 45614
rect 28142 45666 28194 45678
rect 28142 45602 28194 45614
rect 28814 45666 28866 45678
rect 28814 45602 28866 45614
rect 29822 45666 29874 45678
rect 29822 45602 29874 45614
rect 34190 45666 34242 45678
rect 34190 45602 34242 45614
rect 44382 45666 44434 45678
rect 44382 45602 44434 45614
rect 49758 45666 49810 45678
rect 49758 45602 49810 45614
rect 54014 45666 54066 45678
rect 54014 45602 54066 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 4958 45330 5010 45342
rect 4958 45266 5010 45278
rect 10558 45330 10610 45342
rect 10558 45266 10610 45278
rect 13806 45330 13858 45342
rect 13806 45266 13858 45278
rect 16382 45330 16434 45342
rect 16382 45266 16434 45278
rect 17726 45330 17778 45342
rect 17726 45266 17778 45278
rect 23214 45330 23266 45342
rect 23214 45266 23266 45278
rect 26686 45330 26738 45342
rect 26686 45266 26738 45278
rect 40798 45330 40850 45342
rect 40798 45266 40850 45278
rect 2718 45218 2770 45230
rect 2718 45154 2770 45166
rect 7310 45218 7362 45230
rect 7310 45154 7362 45166
rect 9774 45218 9826 45230
rect 9774 45154 9826 45166
rect 14030 45218 14082 45230
rect 28366 45218 28418 45230
rect 20626 45166 20638 45218
rect 20690 45166 20702 45218
rect 14030 45154 14082 45166
rect 28366 45154 28418 45166
rect 30942 45218 30994 45230
rect 30942 45154 30994 45166
rect 42366 45218 42418 45230
rect 50306 45166 50318 45218
rect 50370 45166 50382 45218
rect 53778 45166 53790 45218
rect 53842 45166 53854 45218
rect 42366 45154 42418 45166
rect 9998 45106 10050 45118
rect 9998 45042 10050 45054
rect 10222 45106 10274 45118
rect 10222 45042 10274 45054
rect 10446 45106 10498 45118
rect 25790 45106 25842 45118
rect 19954 45054 19966 45106
rect 20018 45054 20030 45106
rect 10446 45042 10498 45054
rect 25790 45042 25842 45054
rect 26014 45106 26066 45118
rect 26014 45042 26066 45054
rect 26238 45106 26290 45118
rect 30270 45106 30322 45118
rect 31054 45106 31106 45118
rect 28130 45054 28142 45106
rect 28194 45054 28206 45106
rect 30594 45054 30606 45106
rect 30658 45054 30670 45106
rect 26238 45042 26290 45054
rect 30270 45042 30322 45054
rect 31054 45042 31106 45054
rect 31278 45106 31330 45118
rect 42030 45106 42082 45118
rect 35298 45054 35310 45106
rect 35362 45054 35374 45106
rect 41570 45054 41582 45106
rect 41634 45054 41646 45106
rect 43810 45054 43822 45106
rect 43874 45054 43886 45106
rect 49634 45054 49646 45106
rect 49698 45054 49710 45106
rect 52994 45054 53006 45106
rect 53058 45054 53070 45106
rect 31278 45042 31330 45054
rect 42030 45042 42082 45054
rect 26126 44994 26178 45006
rect 38558 44994 38610 45006
rect 13682 44942 13694 44994
rect 13746 44942 13758 44994
rect 22754 44942 22766 44994
rect 22818 44942 22830 44994
rect 35970 44942 35982 44994
rect 36034 44942 36046 44994
rect 38098 44942 38110 44994
rect 38162 44942 38174 44994
rect 26126 44930 26178 44942
rect 38558 44930 38610 44942
rect 41806 44994 41858 45006
rect 41806 44930 41858 44942
rect 42254 44994 42306 45006
rect 47070 44994 47122 45006
rect 56366 44994 56418 45006
rect 44482 44942 44494 44994
rect 44546 44942 44558 44994
rect 46610 44942 46622 44994
rect 46674 44942 46686 44994
rect 52434 44942 52446 44994
rect 52498 44942 52510 44994
rect 55906 44942 55918 44994
rect 55970 44942 55982 44994
rect 42254 44930 42306 44942
rect 47070 44930 47122 44942
rect 56366 44930 56418 44942
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 9774 44546 9826 44558
rect 26910 44546 26962 44558
rect 25442 44494 25454 44546
rect 25506 44494 25518 44546
rect 9774 44482 9826 44494
rect 26910 44482 26962 44494
rect 27134 44546 27186 44558
rect 27134 44482 27186 44494
rect 27246 44546 27298 44558
rect 27246 44482 27298 44494
rect 29710 44546 29762 44558
rect 29710 44482 29762 44494
rect 30718 44546 30770 44558
rect 30718 44482 30770 44494
rect 5854 44434 5906 44446
rect 17166 44434 17218 44446
rect 28926 44434 28978 44446
rect 2594 44382 2606 44434
rect 2658 44382 2670 44434
rect 4722 44382 4734 44434
rect 4786 44382 4798 44434
rect 7186 44382 7198 44434
rect 7250 44382 7262 44434
rect 9314 44382 9326 44434
rect 9378 44382 9390 44434
rect 16594 44382 16606 44434
rect 16658 44382 16670 44434
rect 24658 44382 24670 44434
rect 24722 44382 24734 44434
rect 5854 44370 5906 44382
rect 17166 44370 17218 44382
rect 28926 44370 28978 44382
rect 29934 44434 29986 44446
rect 50878 44434 50930 44446
rect 48514 44382 48526 44434
rect 48578 44382 48590 44434
rect 29934 44370 29986 44382
rect 50878 44370 50930 44382
rect 52670 44434 52722 44446
rect 54674 44382 54686 44434
rect 54738 44382 54750 44434
rect 52670 44370 52722 44382
rect 20862 44322 20914 44334
rect 25902 44322 25954 44334
rect 1922 44270 1934 44322
rect 1986 44270 1998 44322
rect 6402 44270 6414 44322
rect 6466 44270 6478 44322
rect 10098 44270 10110 44322
rect 10162 44270 10174 44322
rect 10322 44270 10334 44322
rect 10386 44270 10398 44322
rect 13794 44270 13806 44322
rect 13858 44270 13870 44322
rect 21746 44270 21758 44322
rect 21810 44270 21822 44322
rect 20862 44258 20914 44270
rect 25902 44258 25954 44270
rect 26014 44322 26066 44334
rect 30830 44322 30882 44334
rect 26226 44270 26238 44322
rect 26290 44270 26302 44322
rect 30146 44270 30158 44322
rect 30210 44270 30222 44322
rect 31042 44270 31054 44322
rect 31106 44270 31118 44322
rect 48066 44270 48078 44322
rect 48130 44270 48142 44322
rect 49074 44270 49086 44322
rect 49138 44270 49150 44322
rect 54002 44270 54014 44322
rect 54066 44270 54078 44322
rect 54450 44270 54462 44322
rect 54514 44270 54526 44322
rect 26014 44258 26066 44270
rect 30830 44258 30882 44270
rect 9886 44210 9938 44222
rect 26798 44210 26850 44222
rect 14466 44158 14478 44210
rect 14530 44158 14542 44210
rect 22530 44158 22542 44210
rect 22594 44158 22606 44210
rect 9886 44146 9938 44158
rect 26798 44146 26850 44158
rect 29598 44210 29650 44222
rect 29598 44146 29650 44158
rect 36206 44210 36258 44222
rect 36206 44146 36258 44158
rect 44606 44210 44658 44222
rect 44606 44146 44658 44158
rect 46398 44210 46450 44222
rect 47394 44158 47406 44210
rect 47458 44158 47470 44210
rect 48962 44158 48974 44210
rect 49026 44158 49038 44210
rect 53442 44158 53454 44210
rect 53506 44158 53518 44210
rect 55122 44158 55134 44210
rect 55186 44158 55198 44210
rect 46398 44146 46450 44158
rect 19294 44098 19346 44110
rect 19294 44034 19346 44046
rect 33966 44098 34018 44110
rect 33966 44034 34018 44046
rect 42366 44098 42418 44110
rect 42366 44034 42418 44046
rect 45838 44098 45890 44110
rect 45838 44034 45890 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 9886 43762 9938 43774
rect 9886 43698 9938 43710
rect 13806 43762 13858 43774
rect 13806 43698 13858 43710
rect 31166 43762 31218 43774
rect 31166 43698 31218 43710
rect 48414 43762 48466 43774
rect 48414 43698 48466 43710
rect 2830 43650 2882 43662
rect 21646 43650 21698 43662
rect 39678 43650 39730 43662
rect 50654 43650 50706 43662
rect 5842 43598 5854 43650
rect 5906 43598 5918 43650
rect 19058 43598 19070 43650
rect 19122 43598 19134 43650
rect 28578 43598 28590 43650
rect 28642 43598 28654 43650
rect 46946 43598 46958 43650
rect 47010 43598 47022 43650
rect 56242 43598 56254 43650
rect 56306 43598 56318 43650
rect 2830 43586 2882 43598
rect 21646 43586 21698 43598
rect 39678 43586 39730 43598
rect 50654 43586 50706 43598
rect 10222 43538 10274 43550
rect 15710 43538 15762 43550
rect 25902 43538 25954 43550
rect 8306 43486 8318 43538
rect 8370 43486 8382 43538
rect 15250 43486 15262 43538
rect 15314 43486 15326 43538
rect 18386 43486 18398 43538
rect 18450 43486 18462 43538
rect 26114 43486 26126 43538
rect 26178 43486 26190 43538
rect 27906 43486 27918 43538
rect 27970 43486 27982 43538
rect 35074 43486 35086 43538
rect 35138 43486 35150 43538
rect 42130 43486 42142 43538
rect 42194 43486 42206 43538
rect 51202 43486 51214 43538
rect 51266 43486 51278 43538
rect 10222 43474 10274 43486
rect 15710 43474 15762 43486
rect 25902 43474 25954 43486
rect 10782 43426 10834 43438
rect 40238 43426 40290 43438
rect 21186 43374 21198 43426
rect 21250 43374 21262 43426
rect 30706 43374 30718 43426
rect 30770 43374 30782 43426
rect 35746 43374 35758 43426
rect 35810 43374 35822 43426
rect 10782 43362 10834 43374
rect 40238 43362 40290 43374
rect 49422 43426 49474 43438
rect 49422 43362 49474 43374
rect 9886 43314 9938 43326
rect 9886 43250 9938 43262
rect 9998 43314 10050 43326
rect 9998 43250 10050 43262
rect 15486 43314 15538 43326
rect 15486 43250 15538 43262
rect 15934 43314 15986 43326
rect 15934 43250 15986 43262
rect 16046 43314 16098 43326
rect 26002 43262 26014 43314
rect 26066 43262 26078 43314
rect 16046 43250 16098 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 14590 42978 14642 42990
rect 9090 42926 9102 42978
rect 9154 42975 9166 42978
rect 9762 42975 9774 42978
rect 9154 42929 9774 42975
rect 9154 42926 9166 42929
rect 9762 42926 9774 42929
rect 9826 42926 9838 42978
rect 14242 42926 14254 42978
rect 14306 42926 14318 42978
rect 14590 42914 14642 42926
rect 18846 42866 18898 42878
rect 42366 42866 42418 42878
rect 52334 42866 52386 42878
rect 2818 42814 2830 42866
rect 2882 42814 2894 42866
rect 4946 42814 4958 42866
rect 5010 42814 5022 42866
rect 8866 42814 8878 42866
rect 8930 42814 8942 42866
rect 12898 42814 12910 42866
rect 12962 42814 12974 42866
rect 15362 42814 15374 42866
rect 15426 42814 15438 42866
rect 23538 42814 23550 42866
rect 23602 42814 23614 42866
rect 34402 42814 34414 42866
rect 34466 42814 34478 42866
rect 36530 42814 36542 42866
rect 36594 42814 36606 42866
rect 39442 42814 39454 42866
rect 39506 42814 39518 42866
rect 41570 42814 41582 42866
rect 41634 42814 41646 42866
rect 46274 42814 46286 42866
rect 46338 42814 46350 42866
rect 48402 42814 48414 42866
rect 48466 42814 48478 42866
rect 48962 42814 48974 42866
rect 49026 42814 49038 42866
rect 51090 42814 51102 42866
rect 51154 42814 51166 42866
rect 18846 42802 18898 42814
rect 42366 42802 42418 42814
rect 52334 42802 52386 42814
rect 14814 42754 14866 42766
rect 42254 42754 42306 42766
rect 2146 42702 2158 42754
rect 2210 42702 2222 42754
rect 6066 42702 6078 42754
rect 6130 42702 6142 42754
rect 9986 42702 9998 42754
rect 10050 42702 10062 42754
rect 18274 42702 18286 42754
rect 18338 42702 18350 42754
rect 26450 42702 26462 42754
rect 26514 42702 26526 42754
rect 33618 42702 33630 42754
rect 33682 42702 33694 42754
rect 38770 42702 38782 42754
rect 38834 42702 38846 42754
rect 14814 42690 14866 42702
rect 42254 42690 42306 42702
rect 42590 42754 42642 42766
rect 42590 42690 42642 42702
rect 42814 42754 42866 42766
rect 42814 42690 42866 42702
rect 44718 42754 44770 42766
rect 45602 42702 45614 42754
rect 45666 42702 45678 42754
rect 51874 42702 51886 42754
rect 51938 42702 51950 42754
rect 44718 42690 44770 42702
rect 6738 42590 6750 42642
rect 6802 42590 6814 42642
rect 10770 42590 10782 42642
rect 10834 42590 10846 42642
rect 17490 42590 17502 42642
rect 17554 42590 17566 42642
rect 25666 42590 25678 42642
rect 25730 42590 25742 42642
rect 9326 42530 9378 42542
rect 9326 42466 9378 42478
rect 13582 42530 13634 42542
rect 13582 42466 13634 42478
rect 20302 42530 20354 42542
rect 20302 42466 20354 42478
rect 20862 42530 20914 42542
rect 20862 42466 20914 42478
rect 37550 42530 37602 42542
rect 37550 42466 37602 42478
rect 38110 42530 38162 42542
rect 38110 42466 38162 42478
rect 42702 42530 42754 42542
rect 42702 42466 42754 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 6862 42194 6914 42206
rect 6862 42130 6914 42142
rect 16494 42194 16546 42206
rect 16494 42130 16546 42142
rect 25790 42194 25842 42206
rect 25790 42130 25842 42142
rect 26574 42194 26626 42206
rect 26574 42130 26626 42142
rect 44942 42194 44994 42206
rect 44942 42130 44994 42142
rect 53342 42194 53394 42206
rect 53342 42130 53394 42142
rect 2718 42082 2770 42094
rect 26014 42082 26066 42094
rect 20178 42030 20190 42082
rect 20242 42030 20254 42082
rect 2718 42018 2770 42030
rect 26014 42018 26066 42030
rect 32622 42082 32674 42094
rect 32622 42018 32674 42030
rect 34302 42082 34354 42094
rect 34302 42018 34354 42030
rect 34750 42082 34802 42094
rect 37202 42030 37214 42082
rect 37266 42030 37278 42082
rect 34750 42018 34802 42030
rect 4398 41970 4450 41982
rect 4398 41906 4450 41918
rect 5182 41970 5234 41982
rect 5182 41906 5234 41918
rect 5406 41970 5458 41982
rect 15822 41970 15874 41982
rect 15026 41918 15038 41970
rect 15090 41918 15102 41970
rect 19394 41918 19406 41970
rect 19458 41918 19470 41970
rect 29250 41918 29262 41970
rect 29314 41918 29326 41970
rect 36530 41918 36542 41970
rect 36594 41918 36606 41970
rect 41570 41918 41582 41970
rect 41634 41918 41646 41970
rect 42354 41918 42366 41970
rect 42418 41918 42430 41970
rect 50082 41918 50094 41970
rect 50146 41918 50158 41970
rect 50754 41918 50766 41970
rect 50818 41918 50830 41970
rect 5406 41906 5458 41918
rect 15822 41906 15874 41918
rect 4958 41858 5010 41870
rect 4958 41794 5010 41806
rect 5630 41858 5682 41870
rect 22766 41858 22818 41870
rect 10322 41806 10334 41858
rect 10386 41806 10398 41858
rect 22306 41806 22318 41858
rect 22370 41806 22382 41858
rect 25666 41806 25678 41858
rect 25730 41806 25742 41858
rect 29922 41806 29934 41858
rect 29986 41806 29998 41858
rect 32050 41806 32062 41858
rect 32114 41806 32126 41858
rect 39330 41806 39342 41858
rect 39394 41806 39406 41858
rect 44482 41806 44494 41858
rect 44546 41806 44558 41858
rect 52882 41806 52894 41858
rect 52946 41806 52958 41858
rect 5630 41794 5682 41806
rect 22766 41794 22818 41806
rect 6078 41746 6130 41758
rect 6078 41682 6130 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 22094 41410 22146 41422
rect 35198 41410 35250 41422
rect 23762 41358 23774 41410
rect 23826 41358 23838 41410
rect 22094 41346 22146 41358
rect 35198 41346 35250 41358
rect 35534 41410 35586 41422
rect 35534 41346 35586 41358
rect 5742 41298 5794 41310
rect 21870 41298 21922 41310
rect 35310 41298 35362 41310
rect 2594 41246 2606 41298
rect 2658 41246 2670 41298
rect 4722 41246 4734 41298
rect 4786 41246 4798 41298
rect 11218 41246 11230 41298
rect 11282 41246 11294 41298
rect 20626 41246 20638 41298
rect 20690 41246 20702 41298
rect 32274 41246 32286 41298
rect 32338 41246 32350 41298
rect 34402 41246 34414 41298
rect 34466 41246 34478 41298
rect 5742 41234 5794 41246
rect 21870 41234 21922 41246
rect 35310 41234 35362 41246
rect 12350 41186 12402 41198
rect 22318 41186 22370 41198
rect 35758 41186 35810 41198
rect 1922 41134 1934 41186
rect 1986 41134 1998 41186
rect 8418 41134 8430 41186
rect 8482 41134 8494 41186
rect 17714 41134 17726 41186
rect 17778 41134 17790 41186
rect 21634 41134 21646 41186
rect 21698 41134 21710 41186
rect 22978 41134 22990 41186
rect 23042 41134 23054 41186
rect 31602 41134 31614 41186
rect 31666 41134 31678 41186
rect 42466 41134 42478 41186
rect 42530 41134 42542 41186
rect 12350 41122 12402 41134
rect 22318 41122 22370 41134
rect 35758 41122 35810 41134
rect 11790 41074 11842 41086
rect 22430 41074 22482 41086
rect 23214 41074 23266 41086
rect 9090 41022 9102 41074
rect 9154 41022 9166 41074
rect 18498 41022 18510 41074
rect 18562 41022 18574 41074
rect 22642 41022 22654 41074
rect 22706 41071 22718 41074
rect 22866 41071 22878 41074
rect 22706 41025 22878 41071
rect 22706 41022 22718 41025
rect 22866 41022 22878 41025
rect 22930 41022 22942 41074
rect 11790 41010 11842 41022
rect 22430 41010 22482 41022
rect 23214 41010 23266 41022
rect 23326 41074 23378 41086
rect 23326 41010 23378 41022
rect 30158 41074 30210 41086
rect 40898 41022 40910 41074
rect 40962 41022 40974 41074
rect 30158 41010 30210 41022
rect 13694 40962 13746 40974
rect 13694 40898 13746 40910
rect 24334 40962 24386 40974
rect 24334 40898 24386 40910
rect 27022 40962 27074 40974
rect 27022 40898 27074 40910
rect 35646 40962 35698 40974
rect 35646 40898 35698 40910
rect 38110 40962 38162 40974
rect 38110 40898 38162 40910
rect 44382 40962 44434 40974
rect 44382 40898 44434 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 9774 40626 9826 40638
rect 9774 40562 9826 40574
rect 11678 40626 11730 40638
rect 11678 40562 11730 40574
rect 18062 40626 18114 40638
rect 18062 40562 18114 40574
rect 36990 40626 37042 40638
rect 36990 40562 37042 40574
rect 54126 40626 54178 40638
rect 54126 40562 54178 40574
rect 5854 40514 5906 40526
rect 13010 40462 13022 40514
rect 13074 40462 13086 40514
rect 29250 40462 29262 40514
rect 29314 40462 29326 40514
rect 34402 40462 34414 40514
rect 34466 40462 34478 40514
rect 38546 40462 38558 40514
rect 38610 40462 38622 40514
rect 5854 40450 5906 40462
rect 19070 40402 19122 40414
rect 25678 40402 25730 40414
rect 12338 40350 12350 40402
rect 12402 40350 12414 40402
rect 21074 40350 21086 40402
rect 21138 40350 21150 40402
rect 19070 40338 19122 40350
rect 25678 40338 25730 40350
rect 26686 40402 26738 40414
rect 49534 40402 49586 40414
rect 27234 40350 27246 40402
rect 27298 40350 27310 40402
rect 33618 40350 33630 40402
rect 33682 40350 33694 40402
rect 37874 40350 37886 40402
rect 37938 40350 37950 40402
rect 46610 40350 46622 40402
rect 46674 40350 46686 40402
rect 50866 40350 50878 40402
rect 50930 40350 50942 40402
rect 26686 40338 26738 40350
rect 49534 40338 49586 40350
rect 8094 40290 8146 40302
rect 15138 40238 15150 40290
rect 15202 40238 15214 40290
rect 23538 40238 23550 40290
rect 23602 40238 23614 40290
rect 36530 40238 36542 40290
rect 36594 40238 36606 40290
rect 40674 40238 40686 40290
rect 40738 40238 40750 40290
rect 43698 40238 43710 40290
rect 43762 40238 43774 40290
rect 45826 40238 45838 40290
rect 45890 40238 45902 40290
rect 51538 40238 51550 40290
rect 51602 40238 51614 40290
rect 53666 40238 53678 40290
rect 53730 40238 53742 40290
rect 8094 40226 8146 40238
rect 49758 40178 49810 40190
rect 50082 40126 50094 40178
rect 50146 40126 50158 40178
rect 49758 40114 49810 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 12462 39730 12514 39742
rect 10434 39678 10446 39730
rect 10498 39678 10510 39730
rect 19954 39678 19966 39730
rect 20018 39678 20030 39730
rect 22978 39678 22990 39730
rect 23042 39678 23054 39730
rect 25106 39678 25118 39730
rect 25170 39678 25182 39730
rect 25666 39678 25678 39730
rect 25730 39678 25742 39730
rect 27794 39678 27806 39730
rect 27858 39678 27870 39730
rect 32498 39678 32510 39730
rect 32562 39678 32574 39730
rect 43810 39678 43822 39730
rect 43874 39678 43886 39730
rect 47618 39678 47630 39730
rect 47682 39678 47694 39730
rect 53666 39678 53678 39730
rect 53730 39678 53742 39730
rect 12462 39666 12514 39678
rect 32958 39618 33010 39630
rect 7634 39566 7646 39618
rect 7698 39566 7710 39618
rect 17154 39566 17166 39618
rect 17218 39566 17230 39618
rect 22306 39566 22318 39618
rect 22370 39566 22382 39618
rect 28578 39566 28590 39618
rect 28642 39566 28654 39618
rect 29698 39566 29710 39618
rect 29762 39566 29774 39618
rect 40898 39566 40910 39618
rect 40962 39566 40974 39618
rect 51202 39566 51214 39618
rect 51266 39566 51278 39618
rect 32958 39554 33010 39566
rect 45614 39506 45666 39518
rect 8306 39454 8318 39506
rect 8370 39454 8382 39506
rect 17826 39454 17838 39506
rect 17890 39454 17902 39506
rect 30370 39454 30382 39506
rect 30434 39454 30446 39506
rect 41682 39454 41694 39506
rect 41746 39454 41758 39506
rect 45614 39442 45666 39454
rect 53454 39506 53506 39518
rect 53454 39442 53506 39454
rect 53678 39506 53730 39518
rect 53678 39442 53730 39454
rect 10894 39394 10946 39406
rect 10894 39330 10946 39342
rect 13806 39394 13858 39406
rect 13806 39330 13858 39342
rect 20862 39394 20914 39406
rect 20862 39330 20914 39342
rect 21534 39394 21586 39406
rect 21534 39330 21586 39342
rect 37662 39394 37714 39406
rect 37662 39330 37714 39342
rect 40014 39394 40066 39406
rect 40014 39330 40066 39342
rect 46846 39394 46898 39406
rect 46846 39330 46898 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 8542 39058 8594 39070
rect 17950 39058 18002 39070
rect 10322 39006 10334 39058
rect 10386 39006 10398 39058
rect 8542 38994 8594 39006
rect 17950 38994 18002 39006
rect 26910 39058 26962 39070
rect 26910 38994 26962 39006
rect 41918 39058 41970 39070
rect 41918 38994 41970 39006
rect 43374 39058 43426 39070
rect 43374 38994 43426 39006
rect 44046 39058 44098 39070
rect 44046 38994 44098 39006
rect 47630 39058 47682 39070
rect 47630 38994 47682 39006
rect 49646 39058 49698 39070
rect 49646 38994 49698 39006
rect 51326 39058 51378 39070
rect 51326 38994 51378 39006
rect 52334 39058 52386 39070
rect 52334 38994 52386 39006
rect 12238 38946 12290 38958
rect 25678 38946 25730 38958
rect 5618 38894 5630 38946
rect 5682 38894 5694 38946
rect 9874 38894 9886 38946
rect 9938 38894 9950 38946
rect 11330 38894 11342 38946
rect 11394 38894 11406 38946
rect 13570 38894 13582 38946
rect 13634 38894 13646 38946
rect 20962 38894 20974 38946
rect 21026 38894 21038 38946
rect 12238 38882 12290 38894
rect 25678 38882 25730 38894
rect 33630 38946 33682 38958
rect 33630 38882 33682 38894
rect 40574 38946 40626 38958
rect 40574 38882 40626 38894
rect 54014 38946 54066 38958
rect 54014 38882 54066 38894
rect 27022 38834 27074 38846
rect 31614 38834 31666 38846
rect 43486 38834 43538 38846
rect 44158 38834 44210 38846
rect 4946 38782 4958 38834
rect 5010 38782 5022 38834
rect 9762 38782 9774 38834
rect 9826 38782 9838 38834
rect 10770 38782 10782 38834
rect 10834 38782 10846 38834
rect 12786 38782 12798 38834
rect 12850 38782 12862 38834
rect 20290 38782 20302 38834
rect 20354 38782 20366 38834
rect 26786 38782 26798 38834
rect 26850 38782 26862 38834
rect 28354 38782 28366 38834
rect 28418 38782 28430 38834
rect 35074 38782 35086 38834
rect 35138 38782 35150 38834
rect 42914 38782 42926 38834
rect 42978 38782 42990 38834
rect 43138 38782 43150 38834
rect 43202 38782 43214 38834
rect 43922 38782 43934 38834
rect 43986 38782 43998 38834
rect 27022 38770 27074 38782
rect 31614 38770 31666 38782
rect 43486 38770 43538 38782
rect 44158 38770 44210 38782
rect 44606 38834 44658 38846
rect 44606 38770 44658 38782
rect 47742 38834 47794 38846
rect 49758 38834 49810 38846
rect 51662 38834 51714 38846
rect 48402 38782 48414 38834
rect 48466 38782 48478 38834
rect 49522 38782 49534 38834
rect 49586 38782 49598 38834
rect 51202 38782 51214 38834
rect 51266 38782 51278 38834
rect 47742 38770 47794 38782
rect 49758 38770 49810 38782
rect 51662 38770 51714 38782
rect 53006 38834 53058 38846
rect 54338 38782 54350 38834
rect 54402 38782 54414 38834
rect 53006 38770 53058 38782
rect 23550 38722 23602 38734
rect 44382 38722 44434 38734
rect 51438 38722 51490 38734
rect 7746 38670 7758 38722
rect 7810 38670 7822 38722
rect 15698 38670 15710 38722
rect 15762 38670 15774 38722
rect 23090 38670 23102 38722
rect 23154 38670 23166 38722
rect 29026 38670 29038 38722
rect 29090 38670 29102 38722
rect 31154 38670 31166 38722
rect 31218 38670 31230 38722
rect 36978 38670 36990 38722
rect 37042 38670 37054 38722
rect 48514 38670 48526 38722
rect 48578 38670 48590 38722
rect 23550 38658 23602 38670
rect 44382 38658 44434 38670
rect 51438 38658 51490 38670
rect 53342 38722 53394 38734
rect 53342 38658 53394 38670
rect 54126 38722 54178 38734
rect 54126 38658 54178 38670
rect 27246 38610 27298 38622
rect 27246 38546 27298 38558
rect 27470 38610 27522 38622
rect 27470 38546 27522 38558
rect 47854 38610 47906 38622
rect 47854 38546 47906 38558
rect 48750 38610 48802 38622
rect 48750 38546 48802 38558
rect 49982 38610 50034 38622
rect 49982 38546 50034 38558
rect 52894 38610 52946 38622
rect 52894 38546 52946 38558
rect 53230 38610 53282 38622
rect 53230 38546 53282 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 15710 38274 15762 38286
rect 52658 38222 52670 38274
rect 52722 38222 52734 38274
rect 15710 38210 15762 38222
rect 12686 38162 12738 38174
rect 36318 38162 36370 38174
rect 25330 38110 25342 38162
rect 25394 38110 25406 38162
rect 27458 38110 27470 38162
rect 27522 38110 27534 38162
rect 32834 38110 32846 38162
rect 32898 38110 32910 38162
rect 34962 38110 34974 38162
rect 35026 38110 35038 38162
rect 12686 38098 12738 38110
rect 36318 38098 36370 38110
rect 36654 38162 36706 38174
rect 52110 38162 52162 38174
rect 37538 38110 37550 38162
rect 37602 38110 37614 38162
rect 39666 38110 39678 38162
rect 39730 38110 39742 38162
rect 41794 38110 41806 38162
rect 41858 38110 41870 38162
rect 43922 38110 43934 38162
rect 43986 38110 43998 38162
rect 47170 38110 47182 38162
rect 47234 38110 47246 38162
rect 49298 38110 49310 38162
rect 49362 38110 49374 38162
rect 54226 38110 54238 38162
rect 54290 38110 54302 38162
rect 56354 38110 56366 38162
rect 56418 38110 56430 38162
rect 36654 38098 36706 38110
rect 52110 38098 52162 38110
rect 15934 38050 15986 38062
rect 8306 37998 8318 38050
rect 8370 37998 8382 38050
rect 15474 37998 15486 38050
rect 15538 37998 15550 38050
rect 15934 37986 15986 37998
rect 16158 38050 16210 38062
rect 36430 38050 36482 38062
rect 50654 38050 50706 38062
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 32162 37998 32174 38050
rect 32226 37998 32238 38050
rect 40338 37998 40350 38050
rect 40402 37998 40414 38050
rect 41010 37998 41022 38050
rect 41074 37998 41086 38050
rect 49970 37998 49982 38050
rect 50034 37998 50046 38050
rect 16158 37986 16210 37998
rect 36430 37986 36482 37998
rect 50654 37986 50706 37998
rect 52334 38050 52386 38062
rect 53442 37998 53454 38050
rect 53506 37998 53518 38050
rect 52334 37986 52386 37998
rect 29598 37938 29650 37950
rect 8978 37886 8990 37938
rect 9042 37886 9054 37938
rect 29598 37874 29650 37886
rect 30382 37938 30434 37950
rect 30382 37874 30434 37886
rect 36766 37938 36818 37950
rect 36766 37874 36818 37886
rect 50990 37938 51042 37950
rect 50990 37874 51042 37886
rect 15598 37826 15650 37838
rect 15598 37762 15650 37774
rect 27918 37826 27970 37838
rect 27918 37762 27970 37774
rect 35534 37826 35586 37838
rect 35534 37762 35586 37774
rect 44606 37826 44658 37838
rect 44606 37762 44658 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 8766 37490 8818 37502
rect 8766 37426 8818 37438
rect 11230 37490 11282 37502
rect 11230 37426 11282 37438
rect 24222 37490 24274 37502
rect 24222 37426 24274 37438
rect 38334 37490 38386 37502
rect 38334 37426 38386 37438
rect 40686 37490 40738 37502
rect 40686 37426 40738 37438
rect 41470 37490 41522 37502
rect 50082 37438 50094 37490
rect 50146 37438 50158 37490
rect 41470 37426 41522 37438
rect 10110 37378 10162 37390
rect 15934 37378 15986 37390
rect 12562 37326 12574 37378
rect 12626 37326 12638 37378
rect 10110 37314 10162 37326
rect 15934 37314 15986 37326
rect 24894 37378 24946 37390
rect 52558 37378 52610 37390
rect 27682 37326 27694 37378
rect 27746 37326 27758 37378
rect 34626 37326 34638 37378
rect 34690 37326 34702 37378
rect 37426 37326 37438 37378
rect 37490 37326 37502 37378
rect 44930 37326 44942 37378
rect 44994 37326 45006 37378
rect 24894 37314 24946 37326
rect 52558 37314 52610 37326
rect 52670 37378 52722 37390
rect 52670 37314 52722 37326
rect 52782 37378 52834 37390
rect 52782 37314 52834 37326
rect 53454 37378 53506 37390
rect 53454 37314 53506 37326
rect 53678 37378 53730 37390
rect 53678 37314 53730 37326
rect 31950 37266 32002 37278
rect 37326 37266 37378 37278
rect 5394 37214 5406 37266
rect 5458 37214 5470 37266
rect 11778 37214 11790 37266
rect 11842 37214 11854 37266
rect 26674 37214 26686 37266
rect 26738 37214 26750 37266
rect 31714 37214 31726 37266
rect 31778 37214 31790 37266
rect 33842 37214 33854 37266
rect 33906 37214 33918 37266
rect 31950 37202 32002 37214
rect 37326 37202 37378 37214
rect 37662 37266 37714 37278
rect 48190 37266 48242 37278
rect 37874 37214 37886 37266
rect 37938 37214 37950 37266
rect 45602 37214 45614 37266
rect 45666 37214 45678 37266
rect 37662 37202 37714 37214
rect 48190 37202 48242 37214
rect 48526 37266 48578 37278
rect 48526 37202 48578 37214
rect 49534 37266 49586 37278
rect 49534 37202 49586 37214
rect 49758 37266 49810 37278
rect 49758 37202 49810 37214
rect 51102 37266 51154 37278
rect 51102 37202 51154 37214
rect 51326 37266 51378 37278
rect 53566 37266 53618 37278
rect 51538 37214 51550 37266
rect 51602 37214 51614 37266
rect 51326 37202 51378 37214
rect 53566 37202 53618 37214
rect 17726 37154 17778 37166
rect 6178 37102 6190 37154
rect 6242 37102 6254 37154
rect 8306 37102 8318 37154
rect 8370 37102 8382 37154
rect 14690 37102 14702 37154
rect 14754 37102 14766 37154
rect 17726 37090 17778 37102
rect 32510 37154 32562 37166
rect 42366 37154 42418 37166
rect 46174 37154 46226 37166
rect 36754 37102 36766 37154
rect 36818 37102 36830 37154
rect 42802 37102 42814 37154
rect 42866 37102 42878 37154
rect 52098 37102 52110 37154
rect 52162 37102 52174 37154
rect 32510 37090 32562 37102
rect 42366 37090 42418 37102
rect 46174 37090 46226 37102
rect 32174 37042 32226 37054
rect 32174 36978 32226 36990
rect 32398 37042 32450 37054
rect 32398 36978 32450 36990
rect 48078 37042 48130 37054
rect 48078 36978 48130 36990
rect 48414 37042 48466 37054
rect 48414 36978 48466 36990
rect 50990 37042 51042 37054
rect 50990 36978 51042 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 7758 36706 7810 36718
rect 7758 36642 7810 36654
rect 8654 36706 8706 36718
rect 8654 36642 8706 36654
rect 7982 36594 8034 36606
rect 27918 36594 27970 36606
rect 9090 36542 9102 36594
rect 9154 36542 9166 36594
rect 11218 36542 11230 36594
rect 11282 36542 11294 36594
rect 15250 36542 15262 36594
rect 15314 36542 15326 36594
rect 17378 36542 17390 36594
rect 17442 36542 17454 36594
rect 20850 36542 20862 36594
rect 20914 36542 20926 36594
rect 25330 36542 25342 36594
rect 25394 36542 25406 36594
rect 27458 36542 27470 36594
rect 27522 36542 27534 36594
rect 7982 36530 8034 36542
rect 27918 36530 27970 36542
rect 35310 36594 35362 36606
rect 35310 36530 35362 36542
rect 37550 36594 37602 36606
rect 42242 36542 42254 36594
rect 42306 36542 42318 36594
rect 48962 36542 48974 36594
rect 49026 36542 49038 36594
rect 50530 36542 50542 36594
rect 50594 36542 50606 36594
rect 52658 36542 52670 36594
rect 52722 36542 52734 36594
rect 37550 36530 37602 36542
rect 8206 36482 8258 36494
rect 12462 36482 12514 36494
rect 43150 36482 43202 36494
rect 12002 36430 12014 36482
rect 12066 36430 12078 36482
rect 14466 36430 14478 36482
rect 14530 36430 14542 36482
rect 17938 36430 17950 36482
rect 18002 36430 18014 36482
rect 24546 36430 24558 36482
rect 24610 36430 24622 36482
rect 39442 36430 39454 36482
rect 39506 36430 39518 36482
rect 42914 36430 42926 36482
rect 42978 36430 42990 36482
rect 8206 36418 8258 36430
rect 12462 36418 12514 36430
rect 43150 36418 43202 36430
rect 43374 36482 43426 36494
rect 43374 36418 43426 36430
rect 43598 36482 43650 36494
rect 46050 36430 46062 36482
rect 46114 36430 46126 36482
rect 49858 36430 49870 36482
rect 49922 36430 49934 36482
rect 43598 36418 43650 36430
rect 6414 36370 6466 36382
rect 6414 36306 6466 36318
rect 7534 36370 7586 36382
rect 18722 36318 18734 36370
rect 18786 36318 18798 36370
rect 40114 36318 40126 36370
rect 40178 36318 40190 36370
rect 46834 36318 46846 36370
rect 46898 36318 46910 36370
rect 7534 36306 7586 36318
rect 5742 36258 5794 36270
rect 5742 36194 5794 36206
rect 13918 36258 13970 36270
rect 13918 36194 13970 36206
rect 21982 36258 22034 36270
rect 21982 36194 22034 36206
rect 29598 36258 29650 36270
rect 29598 36194 29650 36206
rect 43038 36258 43090 36270
rect 43038 36194 43090 36206
rect 44270 36258 44322 36270
rect 44270 36194 44322 36206
rect 45502 36258 45554 36270
rect 45502 36194 45554 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 19742 35922 19794 35934
rect 19742 35858 19794 35870
rect 40350 35922 40402 35934
rect 40350 35858 40402 35870
rect 41470 35922 41522 35934
rect 41470 35858 41522 35870
rect 18846 35810 18898 35822
rect 14018 35758 14030 35810
rect 14082 35758 14094 35810
rect 21858 35758 21870 35810
rect 21922 35758 21934 35810
rect 29362 35758 29374 35810
rect 29426 35758 29438 35810
rect 18846 35746 18898 35758
rect 7758 35698 7810 35710
rect 16606 35698 16658 35710
rect 4498 35646 4510 35698
rect 4562 35646 4574 35698
rect 13234 35646 13246 35698
rect 13298 35646 13310 35698
rect 7758 35634 7810 35646
rect 16606 35634 16658 35646
rect 17614 35698 17666 35710
rect 24446 35698 24498 35710
rect 31950 35698 32002 35710
rect 21186 35646 21198 35698
rect 21250 35646 21262 35698
rect 28578 35646 28590 35698
rect 28642 35646 28654 35698
rect 43474 35646 43486 35698
rect 43538 35646 43550 35698
rect 17614 35634 17666 35646
rect 24446 35634 24498 35646
rect 31950 35634 32002 35646
rect 36094 35586 36146 35598
rect 48078 35586 48130 35598
rect 5170 35534 5182 35586
rect 5234 35534 5246 35586
rect 7298 35534 7310 35586
rect 7362 35534 7374 35586
rect 16146 35534 16158 35586
rect 16210 35534 16222 35586
rect 23986 35534 23998 35586
rect 24050 35534 24062 35586
rect 31490 35534 31502 35586
rect 31554 35534 31566 35586
rect 45378 35534 45390 35586
rect 45442 35534 45454 35586
rect 36094 35522 36146 35534
rect 48078 35522 48130 35534
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 22430 35138 22482 35150
rect 22430 35074 22482 35086
rect 22990 35138 23042 35150
rect 22990 35074 23042 35086
rect 23102 35138 23154 35150
rect 23102 35074 23154 35086
rect 13694 35026 13746 35038
rect 16818 34974 16830 35026
rect 16882 34974 16894 35026
rect 35858 34974 35870 35026
rect 35922 34974 35934 35026
rect 40786 34974 40798 35026
rect 40850 34974 40862 35026
rect 41794 34974 41806 35026
rect 41858 34974 41870 35026
rect 43922 34974 43934 35026
rect 43986 34974 43998 35026
rect 48962 34974 48974 35026
rect 49026 34974 49038 35026
rect 13694 34962 13746 34974
rect 22542 34914 22594 34926
rect 14242 34862 14254 34914
rect 14306 34862 14318 34914
rect 22542 34850 22594 34862
rect 22766 34914 22818 34926
rect 33058 34862 33070 34914
rect 33122 34862 33134 34914
rect 37986 34862 37998 34914
rect 38050 34862 38062 34914
rect 44706 34862 44718 34914
rect 44770 34862 44782 34914
rect 46050 34862 46062 34914
rect 46114 34862 46126 34914
rect 22766 34850 22818 34862
rect 33730 34750 33742 34802
rect 33794 34750 33806 34802
rect 38658 34750 38670 34802
rect 38722 34750 38734 34802
rect 46834 34750 46846 34802
rect 46898 34750 46910 34802
rect 24670 34690 24722 34702
rect 24670 34626 24722 34638
rect 30158 34690 30210 34702
rect 30158 34626 30210 34638
rect 36542 34690 36594 34702
rect 36542 34626 36594 34638
rect 41358 34690 41410 34702
rect 41358 34626 41410 34638
rect 45390 34690 45442 34702
rect 45390 34626 45442 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 18286 34354 18338 34366
rect 18286 34290 18338 34302
rect 32622 34354 32674 34366
rect 32622 34290 32674 34302
rect 33854 34354 33906 34366
rect 33854 34290 33906 34302
rect 38894 34354 38946 34366
rect 38894 34290 38946 34302
rect 39454 34354 39506 34366
rect 39454 34290 39506 34302
rect 47742 34354 47794 34366
rect 47742 34290 47794 34302
rect 17726 34242 17778 34254
rect 40798 34242 40850 34254
rect 13682 34190 13694 34242
rect 13746 34190 13758 34242
rect 30034 34190 30046 34242
rect 30098 34190 30110 34242
rect 37426 34190 37438 34242
rect 37490 34190 37502 34242
rect 17726 34178 17778 34190
rect 40798 34178 40850 34190
rect 18734 34130 18786 34142
rect 6178 34078 6190 34130
rect 6242 34078 6254 34130
rect 16706 34078 16718 34130
rect 16770 34078 16782 34130
rect 19618 34078 19630 34130
rect 19682 34078 19694 34130
rect 29362 34078 29374 34130
rect 29426 34078 29438 34130
rect 38210 34078 38222 34130
rect 38274 34078 38286 34130
rect 41906 34078 41918 34130
rect 41970 34078 41982 34130
rect 18734 34066 18786 34078
rect 9774 34018 9826 34030
rect 22990 34018 23042 34030
rect 6850 33966 6862 34018
rect 6914 33966 6926 34018
rect 8978 33966 8990 34018
rect 9042 33966 9054 34018
rect 20402 33966 20414 34018
rect 20466 33966 20478 34018
rect 22530 33966 22542 34018
rect 22594 33966 22606 34018
rect 32162 33966 32174 34018
rect 32226 33966 32238 34018
rect 35298 33966 35310 34018
rect 35362 33966 35374 34018
rect 45378 33966 45390 34018
rect 45442 33966 45454 34018
rect 9774 33954 9826 33966
rect 22990 33954 23042 33966
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 27806 33458 27858 33470
rect 14354 33406 14366 33458
rect 14418 33406 14430 33458
rect 16482 33406 16494 33458
rect 16546 33406 16558 33458
rect 18610 33406 18622 33458
rect 18674 33406 18686 33458
rect 20738 33406 20750 33458
rect 20802 33406 20814 33458
rect 24434 33406 24446 33458
rect 24498 33406 24510 33458
rect 26562 33406 26574 33458
rect 26626 33406 26638 33458
rect 32610 33406 32622 33458
rect 32674 33406 32686 33458
rect 41234 33406 41246 33458
rect 41298 33406 41310 33458
rect 43362 33406 43374 33458
rect 43426 33406 43438 33458
rect 27806 33394 27858 33406
rect 17154 33294 17166 33346
rect 17218 33294 17230 33346
rect 17826 33294 17838 33346
rect 17890 33294 17902 33346
rect 23762 33294 23774 33346
rect 23826 33294 23838 33346
rect 36306 33294 36318 33346
rect 36370 33294 36382 33346
rect 40562 33294 40574 33346
rect 40626 33294 40638 33346
rect 7086 33234 7138 33246
rect 7086 33170 7138 33182
rect 21646 33234 21698 33246
rect 21646 33170 21698 33182
rect 11230 33122 11282 33134
rect 11230 33058 11282 33070
rect 13694 33122 13746 33134
rect 13694 33058 13746 33070
rect 22990 33122 23042 33134
rect 22990 33058 23042 33070
rect 27246 33122 27298 33134
rect 27246 33058 27298 33070
rect 36766 33122 36818 33134
rect 36766 33058 36818 33070
rect 43822 33122 43874 33134
rect 43822 33058 43874 33070
rect 45726 33122 45778 33134
rect 45726 33058 45778 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 12238 32786 12290 32798
rect 12238 32722 12290 32734
rect 16158 32786 16210 32798
rect 16158 32722 16210 32734
rect 29598 32786 29650 32798
rect 29598 32722 29650 32734
rect 33630 32674 33682 32686
rect 13570 32622 13582 32674
rect 13634 32622 13646 32674
rect 22754 32622 22766 32674
rect 22818 32622 22830 32674
rect 28354 32622 28366 32674
rect 28418 32622 28430 32674
rect 33630 32610 33682 32622
rect 36542 32674 36594 32686
rect 36542 32610 36594 32622
rect 37998 32674 38050 32686
rect 37998 32610 38050 32622
rect 46846 32674 46898 32686
rect 46846 32610 46898 32622
rect 49870 32674 49922 32686
rect 49870 32610 49922 32622
rect 21086 32562 21138 32574
rect 35870 32562 35922 32574
rect 12898 32510 12910 32562
rect 12962 32510 12974 32562
rect 17826 32510 17838 32562
rect 17890 32510 17902 32562
rect 22082 32510 22094 32562
rect 22146 32510 22158 32562
rect 29138 32510 29150 32562
rect 29202 32510 29214 32562
rect 21086 32498 21138 32510
rect 35870 32498 35922 32510
rect 36430 32562 36482 32574
rect 42802 32510 42814 32562
rect 42866 32510 42878 32562
rect 36430 32498 36482 32510
rect 46174 32450 46226 32462
rect 15698 32398 15710 32450
rect 15762 32398 15774 32450
rect 18498 32398 18510 32450
rect 18562 32398 18574 32450
rect 20626 32398 20638 32450
rect 20690 32398 20702 32450
rect 24882 32398 24894 32450
rect 24946 32398 24958 32450
rect 26226 32398 26238 32450
rect 26290 32398 26302 32450
rect 43586 32398 43598 32450
rect 43650 32398 43662 32450
rect 45714 32398 45726 32450
rect 45778 32398 45790 32450
rect 46174 32386 46226 32398
rect 35982 32338 36034 32350
rect 35982 32274 36034 32286
rect 36206 32338 36258 32350
rect 36206 32274 36258 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 17166 31890 17218 31902
rect 10770 31838 10782 31890
rect 10834 31838 10846 31890
rect 12898 31838 12910 31890
rect 12962 31838 12974 31890
rect 16594 31838 16606 31890
rect 16658 31838 16670 31890
rect 17166 31826 17218 31838
rect 19406 31890 19458 31902
rect 19406 31826 19458 31838
rect 20862 31890 20914 31902
rect 26898 31838 26910 31890
rect 26962 31838 26974 31890
rect 34738 31838 34750 31890
rect 34802 31838 34814 31890
rect 38322 31838 38334 31890
rect 38386 31838 38398 31890
rect 40450 31838 40462 31890
rect 40514 31838 40526 31890
rect 20862 31826 20914 31838
rect 46846 31778 46898 31790
rect 10098 31726 10110 31778
rect 10162 31726 10174 31778
rect 13794 31726 13806 31778
rect 13858 31726 13870 31778
rect 24098 31726 24110 31778
rect 24162 31726 24174 31778
rect 31938 31726 31950 31778
rect 32002 31726 32014 31778
rect 32610 31726 32622 31778
rect 32674 31726 32686 31778
rect 37538 31726 37550 31778
rect 37602 31726 37614 31778
rect 51202 31726 51214 31778
rect 51266 31726 51278 31778
rect 46846 31714 46898 31726
rect 18286 31666 18338 31678
rect 43822 31666 43874 31678
rect 14466 31614 14478 31666
rect 14530 31614 14542 31666
rect 24770 31614 24782 31666
rect 24834 31614 24846 31666
rect 49522 31614 49534 31666
rect 49586 31614 49598 31666
rect 18286 31602 18338 31614
rect 43822 31602 43874 31614
rect 20302 31554 20354 31566
rect 20302 31490 20354 31502
rect 21646 31554 21698 31566
rect 21646 31490 21698 31502
rect 27358 31554 27410 31566
rect 27358 31490 27410 31502
rect 35198 31554 35250 31566
rect 35198 31490 35250 31502
rect 36766 31554 36818 31566
rect 36766 31490 36818 31502
rect 40910 31554 40962 31566
rect 40910 31490 40962 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 44942 31218 44994 31230
rect 44942 31154 44994 31166
rect 6414 31106 6466 31118
rect 10098 31054 10110 31106
rect 10162 31054 10174 31106
rect 21634 31054 21646 31106
rect 21698 31054 21710 31106
rect 37874 31054 37886 31106
rect 37938 31054 37950 31106
rect 46610 31054 46622 31106
rect 46674 31054 46686 31106
rect 50306 31054 50318 31106
rect 50370 31054 50382 31106
rect 6414 31042 6466 31054
rect 15710 30994 15762 31006
rect 5954 30942 5966 30994
rect 6018 30942 6030 30994
rect 15026 30942 15038 30994
rect 15090 30942 15102 30994
rect 15710 30930 15762 30942
rect 15934 30994 15986 31006
rect 15934 30930 15986 30942
rect 16158 30994 16210 31006
rect 16158 30930 16210 30942
rect 16270 30994 16322 31006
rect 16270 30930 16322 30942
rect 18510 30994 18562 31006
rect 26350 30994 26402 31006
rect 19058 30942 19070 30994
rect 19122 30942 19134 30994
rect 18510 30930 18562 30942
rect 26350 30930 26402 30942
rect 26798 30994 26850 31006
rect 27010 30942 27022 30994
rect 27074 30942 27086 30994
rect 29698 30942 29710 30994
rect 29762 30942 29774 30994
rect 33730 30942 33742 30994
rect 33794 30942 33806 30994
rect 37090 30942 37102 30994
rect 37154 30942 37166 30994
rect 41570 30942 41582 30994
rect 41634 30942 41646 30994
rect 45938 30942 45950 30994
rect 46002 30942 46014 30994
rect 49522 30942 49534 30994
rect 49586 30942 49598 30994
rect 26798 30930 26850 30942
rect 40462 30882 40514 30894
rect 3042 30830 3054 30882
rect 3106 30830 3118 30882
rect 5170 30830 5182 30882
rect 5234 30830 5246 30882
rect 30370 30830 30382 30882
rect 30434 30830 30446 30882
rect 32498 30830 32510 30882
rect 32562 30830 32574 30882
rect 34402 30830 34414 30882
rect 34466 30830 34478 30882
rect 36530 30830 36542 30882
rect 36594 30830 36606 30882
rect 40002 30830 40014 30882
rect 40066 30830 40078 30882
rect 42354 30830 42366 30882
rect 42418 30830 42430 30882
rect 44482 30830 44494 30882
rect 44546 30830 44558 30882
rect 48738 30830 48750 30882
rect 48802 30830 48814 30882
rect 52434 30830 52446 30882
rect 52498 30830 52510 30882
rect 40462 30818 40514 30830
rect 15598 30770 15650 30782
rect 15598 30706 15650 30718
rect 26238 30770 26290 30782
rect 26238 30706 26290 30718
rect 26574 30770 26626 30782
rect 26574 30706 26626 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 20190 30434 20242 30446
rect 20190 30370 20242 30382
rect 49310 30434 49362 30446
rect 49310 30370 49362 30382
rect 49758 30434 49810 30446
rect 49758 30370 49810 30382
rect 20638 30322 20690 30334
rect 19170 30270 19182 30322
rect 19234 30270 19246 30322
rect 20638 30258 20690 30270
rect 21646 30322 21698 30334
rect 21646 30258 21698 30270
rect 32286 30322 32338 30334
rect 32286 30258 32338 30270
rect 32734 30322 32786 30334
rect 32734 30258 32786 30270
rect 33294 30322 33346 30334
rect 49534 30322 49586 30334
rect 48514 30270 48526 30322
rect 48578 30270 48590 30322
rect 33294 30258 33346 30270
rect 49534 30258 49586 30270
rect 6078 30210 6130 30222
rect 5842 30158 5854 30210
rect 5906 30158 5918 30210
rect 6078 30146 6130 30158
rect 6302 30210 6354 30222
rect 6302 30146 6354 30158
rect 15374 30210 15426 30222
rect 20078 30210 20130 30222
rect 16370 30158 16382 30210
rect 16434 30158 16446 30210
rect 15374 30146 15426 30158
rect 20078 30146 20130 30158
rect 20414 30210 20466 30222
rect 44158 30210 44210 30222
rect 38546 30158 38558 30210
rect 38610 30158 38622 30210
rect 45714 30158 45726 30210
rect 45778 30158 45790 30210
rect 49074 30158 49086 30210
rect 49138 30158 49150 30210
rect 20414 30146 20466 30158
rect 44158 30146 44210 30158
rect 13918 30098 13970 30110
rect 20750 30098 20802 30110
rect 17042 30046 17054 30098
rect 17106 30046 17118 30098
rect 13918 30034 13970 30046
rect 20750 30034 20802 30046
rect 24782 30098 24834 30110
rect 24782 30034 24834 30046
rect 30046 30098 30098 30110
rect 30046 30034 30098 30046
rect 34078 30098 34130 30110
rect 43486 30098 43538 30110
rect 40338 30046 40350 30098
rect 40402 30046 40414 30098
rect 46386 30046 46398 30098
rect 46450 30046 46462 30098
rect 34078 30034 34130 30046
rect 43486 30034 43538 30046
rect 5966 29986 6018 29998
rect 5966 29922 6018 29934
rect 23326 29986 23378 29998
rect 23326 29922 23378 29934
rect 28142 29986 28194 29998
rect 28142 29922 28194 29934
rect 30494 29986 30546 29998
rect 30494 29922 30546 29934
rect 31726 29986 31778 29998
rect 31726 29922 31778 29934
rect 49646 29986 49698 29998
rect 49646 29922 49698 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 9662 29650 9714 29662
rect 9662 29586 9714 29598
rect 13134 29650 13186 29662
rect 13134 29586 13186 29598
rect 17726 29650 17778 29662
rect 17726 29586 17778 29598
rect 40798 29650 40850 29662
rect 40798 29586 40850 29598
rect 46510 29650 46562 29662
rect 46510 29586 46562 29598
rect 5182 29538 5234 29550
rect 5182 29474 5234 29486
rect 5406 29538 5458 29550
rect 5406 29474 5458 29486
rect 11566 29538 11618 29550
rect 11566 29474 11618 29486
rect 16942 29538 16994 29550
rect 19282 29486 19294 29538
rect 19346 29486 19358 29538
rect 22754 29486 22766 29538
rect 22818 29486 22830 29538
rect 27234 29486 27246 29538
rect 27298 29486 27310 29538
rect 30706 29486 30718 29538
rect 30770 29486 30782 29538
rect 16942 29474 16994 29486
rect 36990 29426 37042 29438
rect 8978 29374 8990 29426
rect 9042 29374 9054 29426
rect 18610 29374 18622 29426
rect 18674 29374 18686 29426
rect 21970 29374 21982 29426
rect 22034 29374 22046 29426
rect 26562 29374 26574 29426
rect 26626 29374 26638 29426
rect 29922 29374 29934 29426
rect 29986 29374 29998 29426
rect 33730 29374 33742 29426
rect 33794 29374 33806 29426
rect 36990 29362 37042 29374
rect 39454 29426 39506 29438
rect 39454 29362 39506 29374
rect 39678 29426 39730 29438
rect 45614 29426 45666 29438
rect 41570 29374 41582 29426
rect 41634 29374 41646 29426
rect 45154 29374 45166 29426
rect 45218 29374 45230 29426
rect 39678 29362 39730 29374
rect 45614 29362 45666 29374
rect 49758 29426 49810 29438
rect 49758 29362 49810 29374
rect 39118 29314 39170 29326
rect 45390 29314 45442 29326
rect 5506 29262 5518 29314
rect 5570 29262 5582 29314
rect 6066 29262 6078 29314
rect 6130 29262 6142 29314
rect 8194 29262 8206 29314
rect 8258 29262 8270 29314
rect 21410 29262 21422 29314
rect 21474 29262 21486 29314
rect 24882 29262 24894 29314
rect 24946 29262 24958 29314
rect 29362 29262 29374 29314
rect 29426 29262 29438 29314
rect 32834 29262 32846 29314
rect 32898 29262 32910 29314
rect 34402 29262 34414 29314
rect 34466 29262 34478 29314
rect 36530 29262 36542 29314
rect 36594 29262 36606 29314
rect 42354 29262 42366 29314
rect 42418 29262 42430 29314
rect 44482 29262 44494 29314
rect 44546 29262 44558 29314
rect 39118 29250 39170 29262
rect 45390 29250 45442 29262
rect 45950 29314 46002 29326
rect 45950 29250 46002 29262
rect 49534 29314 49586 29326
rect 49534 29250 49586 29262
rect 39230 29202 39282 29214
rect 39230 29138 39282 29150
rect 39790 29202 39842 29214
rect 39790 29138 39842 29150
rect 45838 29202 45890 29214
rect 50082 29150 50094 29202
rect 50146 29150 50158 29202
rect 45838 29138 45890 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 7534 28866 7586 28878
rect 6514 28814 6526 28866
rect 6578 28814 6590 28866
rect 7534 28802 7586 28814
rect 25902 28866 25954 28878
rect 25902 28802 25954 28814
rect 7422 28754 7474 28766
rect 20078 28754 20130 28766
rect 10770 28702 10782 28754
rect 10834 28702 10846 28754
rect 12898 28702 12910 28754
rect 12962 28702 12974 28754
rect 17378 28702 17390 28754
rect 17442 28702 17454 28754
rect 19506 28702 19518 28754
rect 19570 28702 19582 28754
rect 7422 28690 7474 28702
rect 20078 28690 20130 28702
rect 21758 28754 21810 28766
rect 34962 28702 34974 28754
rect 35026 28702 35038 28754
rect 52658 28702 52670 28754
rect 52722 28702 52734 28754
rect 21758 28690 21810 28702
rect 5966 28642 6018 28654
rect 5966 28578 6018 28590
rect 6190 28642 6242 28654
rect 26126 28642 26178 28654
rect 9986 28590 9998 28642
rect 10050 28590 10062 28642
rect 16706 28590 16718 28642
rect 16770 28590 16782 28642
rect 25666 28590 25678 28642
rect 25730 28590 25742 28642
rect 6190 28578 6242 28590
rect 26126 28578 26178 28590
rect 26350 28642 26402 28654
rect 26350 28578 26402 28590
rect 28254 28642 28306 28654
rect 30258 28590 30270 28642
rect 30322 28590 30334 28642
rect 49746 28590 49758 28642
rect 49810 28590 49822 28642
rect 28254 28578 28306 28590
rect 7310 28530 7362 28542
rect 7310 28466 7362 28478
rect 15710 28530 15762 28542
rect 15710 28466 15762 28478
rect 42254 28530 42306 28542
rect 50530 28478 50542 28530
rect 50594 28478 50606 28530
rect 42254 28466 42306 28478
rect 13806 28418 13858 28430
rect 13806 28354 13858 28366
rect 15150 28418 15202 28430
rect 15150 28354 15202 28366
rect 15262 28418 15314 28430
rect 15262 28354 15314 28366
rect 15486 28418 15538 28430
rect 15486 28354 15538 28366
rect 25118 28418 25170 28430
rect 25118 28354 25170 28366
rect 25790 28418 25842 28430
rect 25790 28354 25842 28366
rect 28814 28418 28866 28430
rect 28814 28354 28866 28366
rect 36318 28418 36370 28430
rect 36318 28354 36370 28366
rect 38894 28418 38946 28430
rect 38894 28354 38946 28366
rect 44270 28418 44322 28430
rect 44270 28354 44322 28366
rect 49310 28418 49362 28430
rect 49310 28354 49362 28366
rect 53342 28418 53394 28430
rect 53342 28354 53394 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 21758 28082 21810 28094
rect 21758 28018 21810 28030
rect 32062 28082 32114 28094
rect 32062 28018 32114 28030
rect 34414 28082 34466 28094
rect 34414 28018 34466 28030
rect 6078 27970 6130 27982
rect 6078 27906 6130 27918
rect 6302 27970 6354 27982
rect 22542 27970 22594 27982
rect 41582 27970 41634 27982
rect 13682 27918 13694 27970
rect 13746 27918 13758 27970
rect 20850 27918 20862 27970
rect 20914 27918 20926 27970
rect 21186 27918 21198 27970
rect 21250 27918 21262 27970
rect 30482 27918 30494 27970
rect 30546 27918 30558 27970
rect 36082 27918 36094 27970
rect 36146 27918 36158 27970
rect 44146 27918 44158 27970
rect 44210 27918 44222 27970
rect 6302 27906 6354 27918
rect 22542 27906 22594 27918
rect 41582 27906 41634 27918
rect 20750 27858 20802 27870
rect 13010 27806 13022 27858
rect 13074 27806 13086 27858
rect 20750 27794 20802 27806
rect 21534 27858 21586 27870
rect 21534 27794 21586 27806
rect 25006 27858 25058 27870
rect 31726 27858 31778 27870
rect 25666 27806 25678 27858
rect 25730 27806 25742 27858
rect 31490 27806 31502 27858
rect 31554 27806 31566 27858
rect 25006 27794 25058 27806
rect 31726 27794 31778 27806
rect 32174 27858 32226 27870
rect 46734 27858 46786 27870
rect 35298 27806 35310 27858
rect 35362 27806 35374 27858
rect 43474 27806 43486 27858
rect 43538 27806 43550 27858
rect 32174 27794 32226 27806
rect 46734 27794 46786 27806
rect 48078 27858 48130 27870
rect 49522 27806 49534 27858
rect 49586 27806 49598 27858
rect 48078 27794 48130 27806
rect 16382 27746 16434 27758
rect 48750 27746 48802 27758
rect 15810 27694 15822 27746
rect 15874 27694 15886 27746
rect 38210 27694 38222 27746
rect 38274 27694 38286 27746
rect 46274 27694 46286 27746
rect 46338 27694 46350 27746
rect 52098 27694 52110 27746
rect 52162 27694 52174 27746
rect 16382 27682 16434 27694
rect 48750 27682 48802 27694
rect 6414 27634 6466 27646
rect 6414 27570 6466 27582
rect 31950 27634 32002 27646
rect 31950 27570 32002 27582
rect 48638 27634 48690 27646
rect 48638 27570 48690 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 6526 27298 6578 27310
rect 6526 27234 6578 27246
rect 14702 27298 14754 27310
rect 14702 27234 14754 27246
rect 15038 27298 15090 27310
rect 15038 27234 15090 27246
rect 6302 27186 6354 27198
rect 6302 27122 6354 27134
rect 8990 27186 9042 27198
rect 8990 27122 9042 27134
rect 9438 27186 9490 27198
rect 14814 27186 14866 27198
rect 52446 27186 52498 27198
rect 10770 27134 10782 27186
rect 10834 27134 10846 27186
rect 12898 27134 12910 27186
rect 12962 27134 12974 27186
rect 25554 27134 25566 27186
rect 25618 27134 25630 27186
rect 27682 27134 27694 27186
rect 27746 27134 27758 27186
rect 32274 27134 32286 27186
rect 32338 27134 32350 27186
rect 38658 27134 38670 27186
rect 38722 27134 38734 27186
rect 40786 27134 40798 27186
rect 40850 27134 40862 27186
rect 49298 27134 49310 27186
rect 49362 27134 49374 27186
rect 56690 27134 56702 27186
rect 56754 27134 56766 27186
rect 9438 27122 9490 27134
rect 14814 27122 14866 27134
rect 52446 27122 52498 27134
rect 8542 27074 8594 27086
rect 15262 27074 15314 27086
rect 41806 27074 41858 27086
rect 50094 27074 50146 27086
rect 10098 27022 10110 27074
rect 10162 27022 10174 27074
rect 24882 27022 24894 27074
rect 24946 27022 24958 27074
rect 35074 27022 35086 27074
rect 35138 27022 35150 27074
rect 37874 27022 37886 27074
rect 37938 27022 37950 27074
rect 46498 27022 46510 27074
rect 46562 27022 46574 27074
rect 49858 27022 49870 27074
rect 49922 27022 49934 27074
rect 8542 27010 8594 27022
rect 15262 27010 15314 27022
rect 41806 27010 41858 27022
rect 50094 27010 50146 27022
rect 50206 27074 50258 27086
rect 50206 27010 50258 27022
rect 51662 27074 51714 27086
rect 53778 27022 53790 27074
rect 53842 27022 53854 27074
rect 51662 27010 51714 27022
rect 13582 26962 13634 26974
rect 13582 26898 13634 26910
rect 20974 26962 21026 26974
rect 20974 26898 21026 26910
rect 28142 26962 28194 26974
rect 41694 26962 41746 26974
rect 34402 26910 34414 26962
rect 34466 26910 34478 26962
rect 28142 26898 28194 26910
rect 41694 26898 41746 26910
rect 41918 26962 41970 26974
rect 51214 26962 51266 26974
rect 47170 26910 47182 26962
rect 47234 26910 47246 26962
rect 41918 26898 41970 26910
rect 51214 26898 51266 26910
rect 51550 26962 51602 26974
rect 51550 26898 51602 26910
rect 52334 26962 52386 26974
rect 54562 26910 54574 26962
rect 54626 26910 54638 26962
rect 52334 26898 52386 26910
rect 8206 26850 8258 26862
rect 6850 26798 6862 26850
rect 6914 26798 6926 26850
rect 8206 26786 8258 26798
rect 15150 26850 15202 26862
rect 15150 26786 15202 26798
rect 18286 26850 18338 26862
rect 18286 26786 18338 26798
rect 23214 26850 23266 26862
rect 51326 26850 51378 26862
rect 42354 26798 42366 26850
rect 42418 26798 42430 26850
rect 50642 26798 50654 26850
rect 50706 26798 50718 26850
rect 23214 26786 23266 26798
rect 51326 26786 51378 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 8878 26514 8930 26526
rect 8878 26450 8930 26462
rect 11454 26514 11506 26526
rect 11454 26450 11506 26462
rect 24894 26514 24946 26526
rect 24894 26450 24946 26462
rect 31838 26514 31890 26526
rect 31838 26450 31890 26462
rect 33742 26514 33794 26526
rect 33742 26450 33794 26462
rect 42142 26514 42194 26526
rect 42142 26450 42194 26462
rect 48414 26514 48466 26526
rect 48414 26450 48466 26462
rect 49758 26514 49810 26526
rect 49758 26450 49810 26462
rect 53230 26514 53282 26526
rect 53230 26450 53282 26462
rect 54014 26514 54066 26526
rect 54014 26450 54066 26462
rect 9998 26402 10050 26414
rect 32398 26402 32450 26414
rect 49870 26402 49922 26414
rect 51326 26402 51378 26414
rect 18498 26350 18510 26402
rect 18562 26350 18574 26402
rect 22306 26350 22318 26402
rect 22370 26350 22382 26402
rect 29250 26350 29262 26402
rect 29314 26350 29326 26402
rect 35746 26350 35758 26402
rect 35810 26350 35822 26402
rect 49970 26350 49982 26402
rect 50034 26350 50046 26402
rect 9998 26338 10050 26350
rect 32398 26338 32450 26350
rect 49870 26338 49922 26350
rect 51326 26338 51378 26350
rect 53678 26402 53730 26414
rect 53678 26338 53730 26350
rect 7310 26290 7362 26302
rect 3378 26238 3390 26290
rect 3442 26238 3454 26290
rect 7310 26226 7362 26238
rect 7534 26290 7586 26302
rect 7534 26226 7586 26238
rect 8542 26290 8594 26302
rect 9886 26290 9938 26302
rect 42254 26290 42306 26302
rect 48078 26290 48130 26302
rect 8978 26238 8990 26290
rect 9042 26238 9054 26290
rect 17826 26238 17838 26290
rect 17890 26238 17902 26290
rect 21634 26238 21646 26290
rect 21698 26238 21710 26290
rect 28578 26238 28590 26290
rect 28642 26238 28654 26290
rect 40226 26238 40238 26290
rect 40290 26238 40302 26290
rect 41570 26238 41582 26290
rect 41634 26238 41646 26290
rect 43586 26238 43598 26290
rect 43650 26238 43662 26290
rect 8542 26226 8594 26238
rect 9886 26226 9938 26238
rect 42254 26226 42306 26238
rect 48078 26226 48130 26238
rect 48414 26290 48466 26302
rect 48414 26226 48466 26238
rect 48750 26290 48802 26302
rect 48750 26226 48802 26238
rect 49534 26290 49586 26302
rect 49534 26226 49586 26238
rect 51438 26290 51490 26302
rect 56130 26238 56142 26290
rect 56194 26238 56206 26290
rect 51438 26226 51490 26238
rect 6862 26178 6914 26190
rect 42030 26178 42082 26190
rect 4162 26126 4174 26178
rect 4226 26126 4238 26178
rect 6290 26126 6302 26178
rect 6354 26126 6366 26178
rect 20626 26126 20638 26178
rect 20690 26126 20702 26178
rect 24434 26126 24446 26178
rect 24498 26126 24510 26178
rect 31378 26126 31390 26178
rect 31442 26126 31454 26178
rect 6862 26114 6914 26126
rect 42030 26114 42082 26126
rect 42814 26178 42866 26190
rect 46846 26178 46898 26190
rect 44258 26126 44270 26178
rect 44322 26126 44334 26178
rect 46386 26126 46398 26178
rect 46450 26126 46462 26178
rect 42814 26114 42866 26126
rect 46846 26114 46898 26126
rect 47518 26178 47570 26190
rect 49858 26126 49870 26178
rect 49922 26126 49934 26178
rect 55346 26126 55358 26178
rect 55410 26126 55422 26178
rect 47518 26114 47570 26126
rect 8766 26066 8818 26078
rect 7858 26014 7870 26066
rect 7922 26014 7934 26066
rect 8766 26002 8818 26014
rect 9774 26066 9826 26078
rect 9774 26002 9826 26014
rect 41806 26066 41858 26078
rect 51326 26066 51378 26078
rect 42578 26014 42590 26066
rect 42642 26063 42654 26066
rect 42914 26063 42926 26066
rect 42642 26017 42926 26063
rect 42642 26014 42654 26017
rect 42914 26014 42926 26017
rect 42978 26014 42990 26066
rect 41806 26002 41858 26014
rect 51326 26002 51378 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 6190 25730 6242 25742
rect 6190 25666 6242 25678
rect 6302 25730 6354 25742
rect 6302 25666 6354 25678
rect 6526 25730 6578 25742
rect 6526 25666 6578 25678
rect 6638 25730 6690 25742
rect 6638 25666 6690 25678
rect 20526 25730 20578 25742
rect 20526 25666 20578 25678
rect 20862 25730 20914 25742
rect 20862 25666 20914 25678
rect 44382 25730 44434 25742
rect 44382 25666 44434 25678
rect 50094 25730 50146 25742
rect 50094 25666 50146 25678
rect 11230 25618 11282 25630
rect 20302 25618 20354 25630
rect 25566 25618 25618 25630
rect 50430 25618 50482 25630
rect 7858 25566 7870 25618
rect 7922 25566 7934 25618
rect 9986 25566 9998 25618
rect 10050 25566 10062 25618
rect 18610 25566 18622 25618
rect 18674 25566 18686 25618
rect 22978 25566 22990 25618
rect 23042 25566 23054 25618
rect 25106 25566 25118 25618
rect 25170 25566 25182 25618
rect 32162 25566 32174 25618
rect 32226 25566 32238 25618
rect 34290 25566 34302 25618
rect 34354 25566 34366 25618
rect 40786 25566 40798 25618
rect 40850 25566 40862 25618
rect 42914 25566 42926 25618
rect 42978 25566 42990 25618
rect 45826 25566 45838 25618
rect 45890 25566 45902 25618
rect 11230 25554 11282 25566
rect 20302 25554 20354 25566
rect 25566 25554 25618 25566
rect 50430 25554 50482 25566
rect 20190 25506 20242 25518
rect 10770 25454 10782 25506
rect 10834 25454 10846 25506
rect 15810 25454 15822 25506
rect 15874 25454 15886 25506
rect 20190 25442 20242 25454
rect 20750 25506 20802 25518
rect 34750 25506 34802 25518
rect 48750 25506 48802 25518
rect 22306 25454 22318 25506
rect 22370 25454 22382 25506
rect 31378 25454 31390 25506
rect 31442 25454 31454 25506
rect 40114 25454 40126 25506
rect 40178 25454 40190 25506
rect 45938 25454 45950 25506
rect 46002 25454 46014 25506
rect 49746 25454 49758 25506
rect 49810 25454 49822 25506
rect 51090 25454 51102 25506
rect 51154 25454 51166 25506
rect 51538 25454 51550 25506
rect 51602 25454 51614 25506
rect 52434 25454 52446 25506
rect 52498 25454 52510 25506
rect 20750 25442 20802 25454
rect 34750 25442 34802 25454
rect 48750 25442 48802 25454
rect 37662 25394 37714 25406
rect 16482 25342 16494 25394
rect 16546 25342 16558 25394
rect 37662 25330 37714 25342
rect 44718 25394 44770 25406
rect 44718 25330 44770 25342
rect 45502 25394 45554 25406
rect 45502 25330 45554 25342
rect 49534 25394 49586 25406
rect 49534 25330 49586 25342
rect 49982 25394 50034 25406
rect 49982 25330 50034 25342
rect 50878 25394 50930 25406
rect 51202 25342 51214 25394
rect 51266 25342 51278 25394
rect 50878 25330 50930 25342
rect 13694 25282 13746 25294
rect 13694 25218 13746 25230
rect 19518 25282 19570 25294
rect 19518 25218 19570 25230
rect 28254 25282 28306 25294
rect 28254 25218 28306 25230
rect 38222 25282 38274 25294
rect 38222 25218 38274 25230
rect 43374 25282 43426 25294
rect 43374 25218 43426 25230
rect 44494 25282 44546 25294
rect 44494 25218 44546 25230
rect 48414 25282 48466 25294
rect 48414 25218 48466 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 17726 24946 17778 24958
rect 17726 24882 17778 24894
rect 44942 24946 44994 24958
rect 44942 24882 44994 24894
rect 48862 24946 48914 24958
rect 48862 24882 48914 24894
rect 6974 24834 7026 24846
rect 25678 24834 25730 24846
rect 39678 24834 39730 24846
rect 14914 24782 14926 24834
rect 14978 24782 14990 24834
rect 19618 24782 19630 24834
rect 19682 24782 19694 24834
rect 28130 24782 28142 24834
rect 28194 24782 28206 24834
rect 36978 24782 36990 24834
rect 37042 24782 37054 24834
rect 6974 24770 7026 24782
rect 25678 24770 25730 24782
rect 39678 24770 39730 24782
rect 45502 24834 45554 24846
rect 45502 24770 45554 24782
rect 49534 24834 49586 24846
rect 49534 24770 49586 24782
rect 49870 24834 49922 24846
rect 49870 24770 49922 24782
rect 7298 24670 7310 24722
rect 7362 24670 7374 24722
rect 13010 24670 13022 24722
rect 13074 24670 13086 24722
rect 18834 24670 18846 24722
rect 18898 24670 18910 24722
rect 27458 24670 27470 24722
rect 27522 24670 27534 24722
rect 36194 24670 36206 24722
rect 36258 24670 36270 24722
rect 45826 24670 45838 24722
rect 45890 24670 45902 24722
rect 51202 24670 51214 24722
rect 51266 24670 51278 24722
rect 55346 24670 55358 24722
rect 55410 24670 55422 24722
rect 7086 24610 7138 24622
rect 7086 24546 7138 24558
rect 18286 24610 18338 24622
rect 22206 24610 22258 24622
rect 45614 24610 45666 24622
rect 51886 24610 51938 24622
rect 55918 24610 55970 24622
rect 21746 24558 21758 24610
rect 21810 24558 21822 24610
rect 30258 24558 30270 24610
rect 30322 24558 30334 24610
rect 39106 24558 39118 24610
rect 39170 24558 39182 24610
rect 51426 24558 51438 24610
rect 51490 24558 51502 24610
rect 52434 24558 52446 24610
rect 52498 24558 52510 24610
rect 54562 24558 54574 24610
rect 54626 24558 54638 24610
rect 18286 24546 18338 24558
rect 22206 24546 22258 24558
rect 45614 24546 45666 24558
rect 51886 24546 51938 24558
rect 55918 24546 55970 24558
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 30046 24162 30098 24174
rect 30046 24098 30098 24110
rect 34414 24162 34466 24174
rect 34414 24098 34466 24110
rect 34638 24162 34690 24174
rect 34638 24098 34690 24110
rect 52334 24162 52386 24174
rect 52334 24098 52386 24110
rect 52670 24162 52722 24174
rect 52670 24098 52722 24110
rect 17054 24050 17106 24062
rect 28030 24050 28082 24062
rect 12226 23998 12238 24050
rect 12290 23998 12302 24050
rect 16594 23998 16606 24050
rect 16658 23998 16670 24050
rect 24658 23998 24670 24050
rect 24722 23998 24734 24050
rect 26786 23998 26798 24050
rect 26850 23998 26862 24050
rect 17054 23986 17106 23998
rect 28030 23986 28082 23998
rect 29710 24050 29762 24062
rect 38322 23998 38334 24050
rect 38386 23998 38398 24050
rect 40450 23998 40462 24050
rect 40514 23998 40526 24050
rect 42578 23998 42590 24050
rect 42642 23998 42654 24050
rect 44706 23998 44718 24050
rect 44770 23998 44782 24050
rect 51314 23998 51326 24050
rect 51378 23998 51390 24050
rect 29710 23986 29762 23998
rect 29822 23938 29874 23950
rect 9426 23886 9438 23938
rect 9490 23886 9502 23938
rect 13682 23886 13694 23938
rect 13746 23886 13758 23938
rect 23986 23886 23998 23938
rect 24050 23886 24062 23938
rect 29822 23874 29874 23886
rect 30270 23938 30322 23950
rect 30270 23874 30322 23886
rect 31390 23938 31442 23950
rect 31390 23874 31442 23886
rect 31726 23938 31778 23950
rect 31726 23874 31778 23886
rect 32174 23938 32226 23950
rect 32174 23874 32226 23886
rect 34302 23938 34354 23950
rect 34302 23874 34354 23886
rect 34862 23938 34914 23950
rect 34862 23874 34914 23886
rect 34974 23938 35026 23950
rect 51662 23938 51714 23950
rect 37538 23886 37550 23938
rect 37602 23886 37614 23938
rect 41794 23886 41806 23938
rect 41858 23886 41870 23938
rect 47058 23886 47070 23938
rect 47122 23886 47134 23938
rect 48290 23886 48302 23938
rect 48354 23886 48366 23938
rect 34974 23874 35026 23886
rect 51662 23874 51714 23886
rect 12910 23826 12962 23838
rect 30382 23826 30434 23838
rect 45614 23826 45666 23838
rect 10098 23774 10110 23826
rect 10162 23774 10174 23826
rect 14466 23774 14478 23826
rect 14530 23774 14542 23826
rect 31490 23774 31502 23826
rect 31554 23774 31566 23826
rect 12910 23762 12962 23774
rect 30382 23762 30434 23774
rect 45614 23762 45666 23774
rect 45726 23826 45778 23838
rect 45726 23762 45778 23774
rect 45838 23826 45890 23838
rect 45838 23762 45890 23774
rect 51102 23826 51154 23838
rect 51102 23762 51154 23774
rect 4622 23714 4674 23726
rect 4622 23650 4674 23662
rect 5742 23714 5794 23726
rect 5742 23650 5794 23662
rect 18958 23714 19010 23726
rect 18958 23650 19010 23662
rect 27358 23714 27410 23726
rect 27358 23650 27410 23662
rect 28478 23714 28530 23726
rect 28478 23650 28530 23662
rect 32398 23714 32450 23726
rect 32398 23650 32450 23662
rect 32846 23714 32898 23726
rect 32846 23650 32898 23662
rect 41022 23714 41074 23726
rect 46846 23714 46898 23726
rect 46274 23662 46286 23714
rect 46338 23662 46350 23714
rect 41022 23650 41074 23662
rect 46846 23650 46898 23662
rect 48078 23714 48130 23726
rect 48078 23650 48130 23662
rect 51326 23714 51378 23726
rect 51326 23650 51378 23662
rect 52558 23714 52610 23726
rect 52558 23650 52610 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 10334 23378 10386 23390
rect 10334 23314 10386 23326
rect 11230 23378 11282 23390
rect 11230 23314 11282 23326
rect 16606 23378 16658 23390
rect 16606 23314 16658 23326
rect 26350 23378 26402 23390
rect 26350 23314 26402 23326
rect 48526 23378 48578 23390
rect 51202 23326 51214 23378
rect 51266 23326 51278 23378
rect 48526 23314 48578 23326
rect 9662 23266 9714 23278
rect 16046 23266 16098 23278
rect 23438 23266 23490 23278
rect 3378 23214 3390 23266
rect 3442 23214 3454 23266
rect 13346 23214 13358 23266
rect 13410 23214 13422 23266
rect 20178 23214 20190 23266
rect 20242 23214 20254 23266
rect 38658 23214 38670 23266
rect 38722 23214 38734 23266
rect 44930 23214 44942 23266
rect 44994 23214 45006 23266
rect 9662 23202 9714 23214
rect 16046 23202 16098 23214
rect 23438 23202 23490 23214
rect 12014 23154 12066 23166
rect 48750 23154 48802 23166
rect 2706 23102 2718 23154
rect 2770 23102 2782 23154
rect 6066 23102 6078 23154
rect 6130 23102 6142 23154
rect 12674 23102 12686 23154
rect 12738 23102 12750 23154
rect 19170 23102 19182 23154
rect 19234 23102 19246 23154
rect 26898 23102 26910 23154
rect 26962 23102 26974 23154
rect 36530 23102 36542 23154
rect 36594 23102 36606 23154
rect 37986 23102 37998 23154
rect 38050 23102 38062 23154
rect 42018 23102 42030 23154
rect 42082 23102 42094 23154
rect 12014 23090 12066 23102
rect 48750 23090 48802 23102
rect 49534 23154 49586 23166
rect 49534 23090 49586 23102
rect 49758 23154 49810 23166
rect 52222 23154 52274 23166
rect 50418 23102 50430 23154
rect 50482 23102 50494 23154
rect 49758 23090 49810 23102
rect 52222 23090 52274 23102
rect 52558 23154 52610 23166
rect 52558 23090 52610 23102
rect 52782 23154 52834 23166
rect 52782 23090 52834 23102
rect 47294 23042 47346 23054
rect 5506 22990 5518 23042
rect 5570 22990 5582 23042
rect 6850 22990 6862 23042
rect 6914 22990 6926 23042
rect 8978 22990 8990 23042
rect 9042 22990 9054 23042
rect 15474 22990 15486 23042
rect 15538 22990 15550 23042
rect 28914 22990 28926 23042
rect 28978 22990 28990 23042
rect 33618 22990 33630 23042
rect 33682 22990 33694 23042
rect 35746 22990 35758 23042
rect 35810 22990 35822 23042
rect 40786 22990 40798 23042
rect 40850 22990 40862 23042
rect 47294 22978 47346 22990
rect 48638 23042 48690 23054
rect 48638 22978 48690 22990
rect 51774 23042 51826 23054
rect 51774 22978 51826 22990
rect 52446 23042 52498 23054
rect 52446 22978 52498 22990
rect 51550 22930 51602 22942
rect 51550 22866 51602 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 12350 22594 12402 22606
rect 12350 22530 12402 22542
rect 12574 22594 12626 22606
rect 12574 22530 12626 22542
rect 41582 22594 41634 22606
rect 41582 22530 41634 22542
rect 41918 22594 41970 22606
rect 41918 22530 41970 22542
rect 47182 22594 47234 22606
rect 47182 22530 47234 22542
rect 47742 22594 47794 22606
rect 47742 22530 47794 22542
rect 51662 22594 51714 22606
rect 51662 22530 51714 22542
rect 13582 22482 13634 22494
rect 35086 22482 35138 22494
rect 1810 22430 1822 22482
rect 1874 22430 1886 22482
rect 3938 22430 3950 22482
rect 4002 22430 4014 22482
rect 8418 22430 8430 22482
rect 8482 22430 8494 22482
rect 15250 22430 15262 22482
rect 15314 22430 15326 22482
rect 17378 22430 17390 22482
rect 17442 22430 17454 22482
rect 18722 22430 18734 22482
rect 18786 22430 18798 22482
rect 20850 22430 20862 22482
rect 20914 22430 20926 22482
rect 24546 22430 24558 22482
rect 24610 22430 24622 22482
rect 26674 22430 26686 22482
rect 26738 22430 26750 22482
rect 28802 22430 28814 22482
rect 28866 22430 28878 22482
rect 31826 22430 31838 22482
rect 31890 22430 31902 22482
rect 33954 22430 33966 22482
rect 34018 22430 34030 22482
rect 38658 22430 38670 22482
rect 38722 22430 38734 22482
rect 40786 22430 40798 22482
rect 40850 22430 40862 22482
rect 13582 22418 13634 22430
rect 35086 22418 35138 22430
rect 12014 22370 12066 22382
rect 4722 22318 4734 22370
rect 4786 22318 4798 22370
rect 6626 22318 6638 22370
rect 6690 22318 6702 22370
rect 12014 22306 12066 22318
rect 12126 22370 12178 22382
rect 41806 22370 41858 22382
rect 14578 22318 14590 22370
rect 14642 22318 14654 22370
rect 17938 22318 17950 22370
rect 18002 22318 18014 22370
rect 21634 22318 21646 22370
rect 21698 22318 21710 22370
rect 26002 22318 26014 22370
rect 26066 22318 26078 22370
rect 31154 22318 31166 22370
rect 31218 22318 31230 22370
rect 37986 22318 37998 22370
rect 38050 22318 38062 22370
rect 41346 22318 41358 22370
rect 41410 22318 41422 22370
rect 12126 22306 12178 22318
rect 41806 22306 41858 22318
rect 46174 22370 46226 22382
rect 46174 22306 46226 22318
rect 46958 22370 47010 22382
rect 46958 22306 47010 22318
rect 47966 22370 48018 22382
rect 47966 22306 48018 22318
rect 48078 22370 48130 22382
rect 48078 22306 48130 22318
rect 51214 22370 51266 22382
rect 51426 22318 51438 22370
rect 51490 22318 51502 22370
rect 51986 22318 51998 22370
rect 52050 22318 52062 22370
rect 51214 22306 51266 22318
rect 12686 22258 12738 22270
rect 34638 22258 34690 22270
rect 46510 22258 46562 22270
rect 22418 22206 22430 22258
rect 22482 22206 22494 22258
rect 46274 22206 46286 22258
rect 46338 22206 46350 22258
rect 12686 22194 12738 22206
rect 34638 22194 34690 22206
rect 46510 22194 46562 22206
rect 47630 22258 47682 22270
rect 47630 22194 47682 22206
rect 42366 22146 42418 22158
rect 42366 22082 42418 22094
rect 51998 22146 52050 22158
rect 51998 22082 52050 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 4958 21810 5010 21822
rect 4958 21746 5010 21758
rect 7310 21810 7362 21822
rect 7310 21746 7362 21758
rect 13134 21810 13186 21822
rect 13134 21746 13186 21758
rect 14142 21810 14194 21822
rect 14142 21746 14194 21758
rect 20862 21810 20914 21822
rect 20862 21746 20914 21758
rect 21310 21810 21362 21822
rect 21310 21746 21362 21758
rect 22318 21810 22370 21822
rect 22318 21746 22370 21758
rect 23998 21810 24050 21822
rect 23998 21746 24050 21758
rect 46062 21810 46114 21822
rect 46062 21746 46114 21758
rect 50878 21810 50930 21822
rect 50878 21746 50930 21758
rect 25678 21698 25730 21710
rect 41470 21698 41522 21710
rect 28354 21646 28366 21698
rect 28418 21646 28430 21698
rect 35634 21646 35646 21698
rect 35698 21646 35710 21698
rect 25678 21634 25730 21646
rect 41470 21634 41522 21646
rect 45614 21698 45666 21710
rect 45614 21634 45666 21646
rect 45838 21698 45890 21710
rect 46386 21646 46398 21698
rect 46450 21695 46462 21698
rect 46834 21695 46846 21698
rect 46450 21649 46846 21695
rect 46450 21646 46462 21649
rect 46834 21646 46846 21649
rect 46898 21646 46910 21698
rect 55346 21646 55358 21698
rect 55410 21646 55422 21698
rect 45838 21634 45890 21646
rect 24110 21586 24162 21598
rect 39342 21586 39394 21598
rect 46286 21586 46338 21598
rect 47070 21586 47122 21598
rect 1810 21534 1822 21586
rect 1874 21534 1886 21586
rect 9874 21534 9886 21586
rect 9938 21534 9950 21586
rect 27682 21534 27694 21586
rect 27746 21534 27758 21586
rect 34962 21534 34974 21586
rect 35026 21534 35038 21586
rect 42130 21534 42142 21586
rect 42194 21534 42206 21586
rect 46834 21534 46846 21586
rect 46898 21534 46910 21586
rect 24110 21522 24162 21534
rect 39342 21522 39394 21534
rect 46286 21522 46338 21534
rect 47070 21522 47122 21534
rect 47294 21586 47346 21598
rect 51426 21534 51438 21586
rect 51490 21534 51502 21586
rect 47294 21522 47346 21534
rect 2482 21422 2494 21474
rect 2546 21422 2558 21474
rect 10546 21422 10558 21474
rect 10610 21422 10622 21474
rect 12674 21422 12686 21474
rect 12738 21422 12750 21474
rect 30482 21422 30494 21474
rect 30546 21422 30558 21474
rect 42914 21422 42926 21474
rect 42978 21422 42990 21474
rect 45042 21422 45054 21474
rect 45106 21422 45118 21474
rect 23998 21362 24050 21374
rect 23998 21298 24050 21310
rect 24334 21362 24386 21374
rect 24334 21298 24386 21310
rect 24558 21362 24610 21374
rect 24558 21298 24610 21310
rect 47406 21362 47458 21374
rect 47406 21298 47458 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 5630 20914 5682 20926
rect 32958 20914 33010 20926
rect 45390 20914 45442 20926
rect 11890 20862 11902 20914
rect 11954 20862 11966 20914
rect 20850 20862 20862 20914
rect 20914 20862 20926 20914
rect 23202 20862 23214 20914
rect 23266 20862 23278 20914
rect 25330 20862 25342 20914
rect 25394 20862 25406 20914
rect 28802 20862 28814 20914
rect 28866 20862 28878 20914
rect 32498 20862 32510 20914
rect 32562 20862 32574 20914
rect 36530 20862 36542 20914
rect 36594 20862 36606 20914
rect 42130 20862 42142 20914
rect 42194 20862 42206 20914
rect 5630 20850 5682 20862
rect 32958 20850 33010 20862
rect 45390 20850 45442 20862
rect 46174 20914 46226 20926
rect 48738 20862 48750 20914
rect 48802 20862 48814 20914
rect 50866 20862 50878 20914
rect 50930 20862 50942 20914
rect 46174 20850 46226 20862
rect 9090 20750 9102 20802
rect 9154 20750 9166 20802
rect 17938 20750 17950 20802
rect 18002 20750 18014 20802
rect 22530 20750 22542 20802
rect 22594 20750 22606 20802
rect 26002 20750 26014 20802
rect 26066 20750 26078 20802
rect 29698 20750 29710 20802
rect 29762 20750 29774 20802
rect 33730 20750 33742 20802
rect 33794 20750 33806 20802
rect 39218 20750 39230 20802
rect 39282 20750 39294 20802
rect 45938 20750 45950 20802
rect 46002 20750 46014 20802
rect 48066 20750 48078 20802
rect 48130 20750 48142 20802
rect 46286 20690 46338 20702
rect 9762 20638 9774 20690
rect 9826 20638 9838 20690
rect 18722 20638 18734 20690
rect 18786 20638 18798 20690
rect 26674 20638 26686 20690
rect 26738 20638 26750 20690
rect 30370 20638 30382 20690
rect 30434 20638 30446 20690
rect 34402 20638 34414 20690
rect 34466 20638 34478 20690
rect 40002 20638 40014 20690
rect 40066 20638 40078 20690
rect 46286 20626 46338 20638
rect 3166 20578 3218 20590
rect 3166 20514 3218 20526
rect 3838 20578 3890 20590
rect 3838 20514 3890 20526
rect 6526 20578 6578 20590
rect 6526 20514 6578 20526
rect 12350 20578 12402 20590
rect 12350 20514 12402 20526
rect 14814 20578 14866 20590
rect 14814 20514 14866 20526
rect 15486 20578 15538 20590
rect 15486 20514 15538 20526
rect 17054 20578 17106 20590
rect 17054 20514 17106 20526
rect 21870 20578 21922 20590
rect 21870 20514 21922 20526
rect 37550 20578 37602 20590
rect 37550 20514 37602 20526
rect 38110 20578 38162 20590
rect 38110 20514 38162 20526
rect 38558 20578 38610 20590
rect 38558 20514 38610 20526
rect 42590 20578 42642 20590
rect 42590 20514 42642 20526
rect 51326 20578 51378 20590
rect 51326 20514 51378 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 9886 20242 9938 20254
rect 9886 20178 9938 20190
rect 10670 20242 10722 20254
rect 10670 20178 10722 20190
rect 19518 20242 19570 20254
rect 19518 20178 19570 20190
rect 20638 20242 20690 20254
rect 20638 20178 20690 20190
rect 27470 20242 27522 20254
rect 27470 20178 27522 20190
rect 29822 20242 29874 20254
rect 29822 20178 29874 20190
rect 34302 20242 34354 20254
rect 40574 20242 40626 20254
rect 38546 20190 38558 20242
rect 38610 20190 38622 20242
rect 34302 20178 34354 20190
rect 40574 20178 40626 20190
rect 50542 20242 50594 20254
rect 50542 20178 50594 20190
rect 54910 20242 54962 20254
rect 54910 20178 54962 20190
rect 8990 20130 9042 20142
rect 31166 20130 31218 20142
rect 43710 20130 43762 20142
rect 49982 20130 50034 20142
rect 2930 20078 2942 20130
rect 2994 20078 3006 20130
rect 6402 20078 6414 20130
rect 6466 20078 6478 20130
rect 14690 20078 14702 20130
rect 14754 20078 14766 20130
rect 21970 20078 21982 20130
rect 22034 20078 22046 20130
rect 35634 20078 35646 20130
rect 35698 20078 35710 20130
rect 38434 20078 38446 20130
rect 38498 20078 38510 20130
rect 39890 20078 39902 20130
rect 39954 20078 39966 20130
rect 47282 20078 47294 20130
rect 47346 20078 47358 20130
rect 53666 20078 53678 20130
rect 53730 20078 53742 20130
rect 8990 20066 9042 20078
rect 31166 20066 31218 20078
rect 43710 20066 43762 20078
rect 49982 20066 50034 20078
rect 18062 20018 18114 20030
rect 30942 20018 30994 20030
rect 2146 19966 2158 20018
rect 2210 19966 2222 20018
rect 5618 19966 5630 20018
rect 5682 19966 5694 20018
rect 14018 19966 14030 20018
rect 14082 19966 14094 20018
rect 18498 19966 18510 20018
rect 18562 19966 18574 20018
rect 21186 19966 21198 20018
rect 21250 19966 21262 20018
rect 34850 19966 34862 20018
rect 34914 19966 34926 20018
rect 38322 19966 38334 20018
rect 38386 19966 38398 20018
rect 39330 19966 39342 20018
rect 39394 19966 39406 20018
rect 48066 19966 48078 20018
rect 48130 19966 48142 20018
rect 54450 19966 54462 20018
rect 54514 19966 54526 20018
rect 18062 19954 18114 19966
rect 30942 19954 30994 19966
rect 18286 19906 18338 19918
rect 24558 19906 24610 19918
rect 5058 19854 5070 19906
rect 5122 19854 5134 19906
rect 8530 19854 8542 19906
rect 8594 19854 8606 19906
rect 16818 19854 16830 19906
rect 16882 19854 16894 19906
rect 24098 19854 24110 19906
rect 24162 19854 24174 19906
rect 18286 19842 18338 19854
rect 24558 19842 24610 19854
rect 25566 19906 25618 19918
rect 48526 19906 48578 19918
rect 31266 19854 31278 19906
rect 31330 19854 31342 19906
rect 37762 19854 37774 19906
rect 37826 19854 37838 19906
rect 45154 19854 45166 19906
rect 45218 19854 45230 19906
rect 51538 19854 51550 19906
rect 51602 19854 51614 19906
rect 25566 19842 25618 19854
rect 48526 19842 48578 19854
rect 17726 19794 17778 19806
rect 17726 19730 17778 19742
rect 17838 19794 17890 19806
rect 17838 19730 17890 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 6302 19458 6354 19470
rect 6302 19394 6354 19406
rect 6526 19458 6578 19470
rect 6526 19394 6578 19406
rect 6750 19458 6802 19470
rect 6750 19394 6802 19406
rect 6078 19346 6130 19358
rect 13582 19346 13634 19358
rect 2818 19294 2830 19346
rect 2882 19294 2894 19346
rect 4946 19294 4958 19346
rect 5010 19294 5022 19346
rect 12562 19294 12574 19346
rect 12626 19294 12638 19346
rect 6078 19282 6130 19294
rect 13582 19282 13634 19294
rect 21534 19346 21586 19358
rect 21534 19282 21586 19294
rect 22990 19346 23042 19358
rect 41358 19346 41410 19358
rect 33506 19294 33518 19346
rect 33570 19294 33582 19346
rect 40898 19294 40910 19346
rect 40962 19294 40974 19346
rect 49634 19294 49646 19346
rect 49698 19294 49710 19346
rect 51762 19294 51774 19346
rect 51826 19294 51838 19346
rect 53442 19294 53454 19346
rect 53506 19294 53518 19346
rect 22990 19282 23042 19294
rect 41358 19282 41410 19294
rect 56814 19234 56866 19246
rect 2146 19182 2158 19234
rect 2210 19182 2222 19234
rect 9650 19182 9662 19234
rect 9714 19182 9726 19234
rect 15586 19182 15598 19234
rect 15650 19182 15662 19234
rect 23538 19182 23550 19234
rect 23602 19182 23614 19234
rect 30594 19182 30606 19234
rect 30658 19182 30670 19234
rect 38098 19182 38110 19234
rect 38162 19182 38174 19234
rect 48850 19182 48862 19234
rect 48914 19182 48926 19234
rect 56242 19182 56254 19234
rect 56306 19182 56318 19234
rect 56814 19170 56866 19182
rect 52670 19122 52722 19134
rect 10434 19070 10446 19122
rect 10498 19070 10510 19122
rect 20066 19070 20078 19122
rect 20130 19070 20142 19122
rect 25554 19070 25566 19122
rect 25618 19070 25630 19122
rect 31378 19070 31390 19122
rect 31442 19070 31454 19122
rect 38770 19070 38782 19122
rect 38834 19070 38846 19122
rect 55570 19070 55582 19122
rect 55634 19070 55646 19122
rect 52670 19058 52722 19070
rect 7198 19010 7250 19022
rect 7198 18946 7250 18958
rect 33966 19010 34018 19022
rect 33966 18946 34018 18958
rect 46510 19010 46562 19022
rect 46510 18946 46562 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 5294 18674 5346 18686
rect 5294 18610 5346 18622
rect 10670 18674 10722 18686
rect 10670 18610 10722 18622
rect 31614 18674 31666 18686
rect 31614 18610 31666 18622
rect 38894 18674 38946 18686
rect 38894 18610 38946 18622
rect 53678 18674 53730 18686
rect 53678 18610 53730 18622
rect 13246 18562 13298 18574
rect 13246 18498 13298 18510
rect 23662 18562 23714 18574
rect 54798 18562 54850 18574
rect 43922 18510 43934 18562
rect 43986 18510 43998 18562
rect 23662 18498 23714 18510
rect 54798 18498 54850 18510
rect 13134 18450 13186 18462
rect 21310 18450 21362 18462
rect 37438 18450 37490 18462
rect 7634 18398 7646 18450
rect 7698 18398 7710 18450
rect 7858 18398 7870 18450
rect 7922 18398 7934 18450
rect 8194 18398 8206 18450
rect 8258 18398 8270 18450
rect 13458 18398 13470 18450
rect 13522 18398 13534 18450
rect 14130 18398 14142 18450
rect 14194 18398 14206 18450
rect 17938 18398 17950 18450
rect 18002 18398 18014 18450
rect 21746 18398 21758 18450
rect 21810 18398 21822 18450
rect 25666 18398 25678 18450
rect 25730 18398 25742 18450
rect 34066 18398 34078 18450
rect 34130 18398 34142 18450
rect 13134 18386 13186 18398
rect 21310 18386 21362 18398
rect 37438 18386 37490 18398
rect 40798 18450 40850 18462
rect 53342 18450 53394 18462
rect 41906 18398 41918 18450
rect 41970 18398 41982 18450
rect 49634 18398 49646 18450
rect 49698 18398 49710 18450
rect 50306 18398 50318 18450
rect 50370 18398 50382 18450
rect 40798 18386 40850 18398
rect 53342 18386 53394 18398
rect 53566 18450 53618 18462
rect 53566 18386 53618 18398
rect 21982 18338 22034 18350
rect 29038 18338 29090 18350
rect 14802 18286 14814 18338
rect 14866 18286 14878 18338
rect 16930 18286 16942 18338
rect 16994 18286 17006 18338
rect 18610 18286 18622 18338
rect 18674 18286 18686 18338
rect 20738 18286 20750 18338
rect 20802 18286 20814 18338
rect 26450 18286 26462 18338
rect 26514 18286 26526 18338
rect 28578 18286 28590 18338
rect 28642 18286 28654 18338
rect 34850 18286 34862 18338
rect 34914 18286 34926 18338
rect 36978 18286 36990 18338
rect 37042 18286 37054 18338
rect 52434 18286 52446 18338
rect 52498 18286 52510 18338
rect 21982 18274 22034 18286
rect 29038 18274 29090 18286
rect 22206 18226 22258 18238
rect 8418 18174 8430 18226
rect 8482 18174 8494 18226
rect 12674 18174 12686 18226
rect 12738 18174 12750 18226
rect 22206 18162 22258 18174
rect 22430 18226 22482 18238
rect 22430 18162 22482 18174
rect 22542 18226 22594 18238
rect 22542 18162 22594 18174
rect 53230 18226 53282 18238
rect 53230 18162 53282 18174
rect 53790 18226 53842 18238
rect 53790 18162 53842 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 13582 17778 13634 17790
rect 12674 17726 12686 17778
rect 12738 17726 12750 17778
rect 13582 17714 13634 17726
rect 17278 17778 17330 17790
rect 57150 17778 57202 17790
rect 22642 17726 22654 17778
rect 22706 17726 22718 17778
rect 24770 17726 24782 17778
rect 24834 17726 24846 17778
rect 44482 17726 44494 17778
rect 44546 17726 44558 17778
rect 45490 17726 45502 17778
rect 45554 17726 45566 17778
rect 47618 17726 47630 17778
rect 47682 17726 47694 17778
rect 53778 17726 53790 17778
rect 53842 17726 53854 17778
rect 55906 17726 55918 17778
rect 55970 17726 55982 17778
rect 17278 17714 17330 17726
rect 57150 17714 57202 17726
rect 8306 17614 8318 17666
rect 8370 17614 8382 17666
rect 25442 17614 25454 17666
rect 25506 17614 25518 17666
rect 41682 17614 41694 17666
rect 41746 17614 41758 17666
rect 48290 17614 48302 17666
rect 48354 17614 48366 17666
rect 56690 17614 56702 17666
rect 56754 17614 56766 17666
rect 18846 17554 18898 17566
rect 18846 17490 18898 17502
rect 26462 17554 26514 17566
rect 26462 17490 26514 17502
rect 35086 17554 35138 17566
rect 35086 17490 35138 17502
rect 41022 17554 41074 17566
rect 42354 17502 42366 17554
rect 42418 17502 42430 17554
rect 41022 17490 41074 17502
rect 6526 17442 6578 17454
rect 6526 17378 6578 17390
rect 20190 17442 20242 17454
rect 20190 17378 20242 17390
rect 29598 17442 29650 17454
rect 29598 17378 29650 17390
rect 48862 17442 48914 17454
rect 48862 17378 48914 17390
rect 51998 17442 52050 17454
rect 51998 17378 52050 17390
rect 52670 17442 52722 17454
rect 52670 17378 52722 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 22654 17106 22706 17118
rect 22654 17042 22706 17054
rect 25790 17106 25842 17118
rect 25790 17042 25842 17054
rect 27582 17106 27634 17118
rect 36766 17106 36818 17118
rect 34738 17054 34750 17106
rect 34802 17054 34814 17106
rect 27582 17042 27634 17054
rect 36766 17042 36818 17054
rect 48750 17106 48802 17118
rect 48750 17042 48802 17054
rect 9774 16994 9826 17006
rect 6402 16942 6414 16994
rect 6466 16942 6478 16994
rect 9774 16930 9826 16942
rect 14926 16994 14978 17006
rect 14926 16930 14978 16942
rect 17726 16994 17778 17006
rect 31614 16994 31666 17006
rect 39790 16994 39842 17006
rect 20066 16942 20078 16994
rect 20130 16942 20142 16994
rect 33730 16942 33742 16994
rect 33794 16942 33806 16994
rect 35186 16942 35198 16994
rect 35250 16942 35262 16994
rect 37314 16942 37326 16994
rect 37378 16942 37390 16994
rect 43474 16942 43486 16994
rect 43538 16942 43550 16994
rect 51538 16942 51550 16994
rect 51602 16942 51614 16994
rect 17726 16930 17778 16942
rect 31614 16930 31666 16942
rect 39790 16930 39842 16942
rect 8990 16882 9042 16894
rect 5058 16830 5070 16882
rect 5122 16830 5134 16882
rect 5730 16830 5742 16882
rect 5794 16830 5806 16882
rect 8990 16818 9042 16830
rect 10782 16882 10834 16894
rect 23326 16882 23378 16894
rect 46062 16882 46114 16894
rect 11442 16830 11454 16882
rect 11506 16830 11518 16882
rect 19394 16830 19406 16882
rect 19458 16830 19470 16882
rect 28130 16830 28142 16882
rect 28194 16830 28206 16882
rect 28914 16830 28926 16882
rect 28978 16830 28990 16882
rect 33618 16830 33630 16882
rect 33682 16830 33694 16882
rect 34626 16830 34638 16882
rect 34690 16830 34702 16882
rect 37538 16830 37550 16882
rect 37602 16830 37614 16882
rect 38210 16830 38222 16882
rect 38274 16830 38286 16882
rect 38546 16830 38558 16882
rect 38610 16830 38622 16882
rect 42802 16830 42814 16882
rect 42866 16830 42878 16882
rect 49522 16830 49534 16882
rect 49586 16830 49598 16882
rect 10782 16818 10834 16830
rect 23326 16818 23378 16830
rect 46062 16818 46114 16830
rect 23550 16770 23602 16782
rect 48302 16770 48354 16782
rect 2146 16718 2158 16770
rect 2210 16718 2222 16770
rect 4274 16718 4286 16770
rect 4338 16718 4350 16770
rect 8530 16718 8542 16770
rect 8594 16718 8606 16770
rect 12114 16718 12126 16770
rect 12178 16718 12190 16770
rect 14242 16718 14254 16770
rect 14306 16718 14318 16770
rect 22194 16718 22206 16770
rect 22258 16718 22270 16770
rect 31042 16718 31054 16770
rect 31106 16718 31118 16770
rect 45602 16718 45614 16770
rect 45666 16718 45678 16770
rect 23550 16706 23602 16718
rect 48302 16706 48354 16718
rect 38558 16658 38610 16670
rect 23874 16606 23886 16658
rect 23938 16606 23950 16658
rect 38558 16594 38610 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 13918 16322 13970 16334
rect 13918 16258 13970 16270
rect 14142 16322 14194 16334
rect 14142 16258 14194 16270
rect 37662 16322 37714 16334
rect 37662 16258 37714 16270
rect 37998 16322 38050 16334
rect 37998 16258 38050 16270
rect 5630 16210 5682 16222
rect 12798 16210 12850 16222
rect 9426 16158 9438 16210
rect 9490 16158 9502 16210
rect 11554 16158 11566 16210
rect 11618 16158 11630 16210
rect 5630 16146 5682 16158
rect 12798 16146 12850 16158
rect 13806 16210 13858 16222
rect 19854 16210 19906 16222
rect 37774 16210 37826 16222
rect 17266 16158 17278 16210
rect 17330 16158 17342 16210
rect 19394 16158 19406 16210
rect 19458 16158 19470 16210
rect 30818 16158 30830 16210
rect 30882 16158 30894 16210
rect 32946 16158 32958 16210
rect 33010 16158 33022 16210
rect 38770 16158 38782 16210
rect 38834 16158 38846 16210
rect 40898 16158 40910 16210
rect 40962 16158 40974 16210
rect 45490 16158 45502 16210
rect 45554 16158 45566 16210
rect 52658 16158 52670 16210
rect 52722 16158 52734 16210
rect 13806 16146 13858 16158
rect 19854 16146 19906 16158
rect 37774 16146 37826 16158
rect 14366 16098 14418 16110
rect 8754 16046 8766 16098
rect 8818 16046 8830 16098
rect 16594 16046 16606 16098
rect 16658 16046 16670 16098
rect 30034 16046 30046 16098
rect 30098 16046 30110 16098
rect 38210 16046 38222 16098
rect 38274 16046 38286 16098
rect 41682 16046 41694 16098
rect 41746 16046 41758 16098
rect 48290 16046 48302 16098
rect 48354 16046 48366 16098
rect 49746 16046 49758 16098
rect 49810 16046 49822 16098
rect 14366 16034 14418 16046
rect 4510 15986 4562 15998
rect 4510 15922 4562 15934
rect 12238 15986 12290 15998
rect 12238 15922 12290 15934
rect 44046 15986 44098 15998
rect 53454 15986 53506 15998
rect 47618 15934 47630 15986
rect 47682 15934 47694 15986
rect 50530 15934 50542 15986
rect 50594 15934 50606 15986
rect 44046 15922 44098 15934
rect 53454 15922 53506 15934
rect 13806 15874 13858 15886
rect 13806 15810 13858 15822
rect 23774 15874 23826 15886
rect 23774 15810 23826 15822
rect 27134 15874 27186 15886
rect 27134 15810 27186 15822
rect 33518 15874 33570 15886
rect 33518 15810 33570 15822
rect 34078 15874 34130 15886
rect 34078 15810 34130 15822
rect 36430 15874 36482 15886
rect 36430 15810 36482 15822
rect 42142 15874 42194 15886
rect 42142 15810 42194 15822
rect 44718 15874 44770 15886
rect 44718 15810 44770 15822
rect 49198 15874 49250 15886
rect 49198 15810 49250 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 38894 15538 38946 15550
rect 38894 15474 38946 15486
rect 52894 15538 52946 15550
rect 52894 15474 52946 15486
rect 53342 15538 53394 15550
rect 53342 15474 53394 15486
rect 42254 15426 42306 15438
rect 15250 15374 15262 15426
rect 15314 15374 15326 15426
rect 26898 15374 26910 15426
rect 26962 15374 26974 15426
rect 36306 15374 36318 15426
rect 36370 15374 36382 15426
rect 42254 15362 42306 15374
rect 48414 15426 48466 15438
rect 54126 15426 54178 15438
rect 50306 15374 50318 15426
rect 50370 15374 50382 15426
rect 48414 15362 48466 15374
rect 54126 15362 54178 15374
rect 18846 15314 18898 15326
rect 45838 15314 45890 15326
rect 16034 15262 16046 15314
rect 16098 15262 16110 15314
rect 19506 15262 19518 15314
rect 19570 15262 19582 15314
rect 26226 15262 26238 15314
rect 26290 15262 26302 15314
rect 35634 15262 35646 15314
rect 35698 15262 35710 15314
rect 45602 15262 45614 15314
rect 45666 15262 45678 15314
rect 18846 15250 18898 15262
rect 45838 15250 45890 15262
rect 46062 15314 46114 15326
rect 46062 15250 46114 15262
rect 46286 15314 46338 15326
rect 49634 15262 49646 15314
rect 49698 15262 49710 15314
rect 46286 15250 46338 15262
rect 10110 15202 10162 15214
rect 16606 15202 16658 15214
rect 13122 15150 13134 15202
rect 13186 15150 13198 15202
rect 21522 15150 21534 15202
rect 21586 15150 21598 15202
rect 29026 15150 29038 15202
rect 29090 15150 29102 15202
rect 38434 15150 38446 15202
rect 38498 15150 38510 15202
rect 52434 15150 52446 15202
rect 52498 15150 52510 15202
rect 10110 15138 10162 15150
rect 16606 15138 16658 15150
rect 9998 15090 10050 15102
rect 9998 15026 10050 15038
rect 46398 15090 46450 15102
rect 52658 15038 52670 15090
rect 52722 15087 52734 15090
rect 53330 15087 53342 15090
rect 52722 15041 53342 15087
rect 52722 15038 52734 15041
rect 53330 15038 53342 15041
rect 53394 15038 53406 15090
rect 46398 15026 46450 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 11342 14642 11394 14654
rect 20190 14642 20242 14654
rect 43822 14642 43874 14654
rect 50766 14642 50818 14654
rect 10770 14590 10782 14642
rect 10834 14590 10846 14642
rect 19730 14590 19742 14642
rect 19794 14590 19806 14642
rect 22530 14590 22542 14642
rect 22594 14590 22606 14642
rect 24658 14590 24670 14642
rect 24722 14590 24734 14642
rect 28130 14590 28142 14642
rect 28194 14590 28206 14642
rect 32722 14590 32734 14642
rect 32786 14590 32798 14642
rect 34850 14590 34862 14642
rect 34914 14590 34926 14642
rect 41682 14590 41694 14642
rect 41746 14590 41758 14642
rect 48178 14590 48190 14642
rect 48242 14590 48254 14642
rect 50306 14590 50318 14642
rect 50370 14590 50382 14642
rect 53442 14590 53454 14642
rect 53506 14590 53518 14642
rect 55570 14590 55582 14642
rect 55634 14590 55646 14642
rect 11342 14578 11394 14590
rect 20190 14578 20242 14590
rect 43822 14578 43874 14590
rect 50766 14578 50818 14590
rect 56814 14530 56866 14542
rect 7970 14478 7982 14530
rect 8034 14478 8046 14530
rect 16818 14478 16830 14530
rect 16882 14478 16894 14530
rect 21746 14478 21758 14530
rect 21810 14478 21822 14530
rect 25330 14478 25342 14530
rect 25394 14478 25406 14530
rect 32050 14478 32062 14530
rect 32114 14478 32126 14530
rect 39554 14478 39566 14530
rect 39618 14478 39630 14530
rect 47506 14478 47518 14530
rect 47570 14478 47582 14530
rect 56354 14478 56366 14530
rect 56418 14478 56430 14530
rect 56814 14466 56866 14478
rect 8642 14366 8654 14418
rect 8706 14366 8718 14418
rect 17602 14366 17614 14418
rect 17666 14366 17678 14418
rect 26002 14366 26014 14418
rect 26066 14366 26078 14418
rect 16270 14306 16322 14318
rect 16270 14242 16322 14254
rect 20862 14306 20914 14318
rect 20862 14242 20914 14254
rect 30046 14306 30098 14318
rect 30046 14242 30098 14254
rect 30942 14306 30994 14318
rect 30942 14242 30994 14254
rect 35310 14306 35362 14318
rect 35310 14242 35362 14254
rect 36318 14306 36370 14318
rect 36318 14242 36370 14254
rect 46286 14306 46338 14318
rect 46286 14242 46338 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 17838 13970 17890 13982
rect 17838 13906 17890 13918
rect 23886 13970 23938 13982
rect 23886 13906 23938 13918
rect 26014 13970 26066 13982
rect 26014 13906 26066 13918
rect 33518 13970 33570 13982
rect 33518 13906 33570 13918
rect 38782 13970 38834 13982
rect 38782 13906 38834 13918
rect 53678 13970 53730 13982
rect 53678 13906 53730 13918
rect 6974 13858 7026 13870
rect 40014 13858 40066 13870
rect 8082 13806 8094 13858
rect 8146 13806 8158 13858
rect 8642 13806 8654 13858
rect 8706 13806 8718 13858
rect 21298 13806 21310 13858
rect 21362 13806 21374 13858
rect 36194 13806 36206 13858
rect 36258 13806 36270 13858
rect 6974 13794 7026 13806
rect 40014 13794 40066 13806
rect 10446 13746 10498 13758
rect 47854 13746 47906 13758
rect 53342 13746 53394 13758
rect 3490 13694 3502 13746
rect 3554 13694 3566 13746
rect 8978 13694 8990 13746
rect 9042 13694 9054 13746
rect 9986 13694 9998 13746
rect 10050 13694 10062 13746
rect 10882 13694 10894 13746
rect 10946 13694 10958 13746
rect 14018 13694 14030 13746
rect 14082 13694 14094 13746
rect 20626 13694 20638 13746
rect 20690 13694 20702 13746
rect 26898 13694 26910 13746
rect 26962 13694 26974 13746
rect 35522 13694 35534 13746
rect 35586 13694 35598 13746
rect 46946 13694 46958 13746
rect 47010 13694 47022 13746
rect 53106 13694 53118 13746
rect 53170 13694 53182 13746
rect 10446 13682 10498 13694
rect 47854 13682 47906 13694
rect 53342 13682 53394 13694
rect 53566 13746 53618 13758
rect 53566 13682 53618 13694
rect 53790 13746 53842 13758
rect 53790 13682 53842 13694
rect 6862 13634 6914 13646
rect 4162 13582 4174 13634
rect 4226 13582 4238 13634
rect 6290 13582 6302 13634
rect 6354 13582 6366 13634
rect 6862 13570 6914 13582
rect 7758 13634 7810 13646
rect 10210 13582 10222 13634
rect 10274 13582 10286 13634
rect 11106 13582 11118 13634
rect 11170 13582 11182 13634
rect 14802 13582 14814 13634
rect 14866 13582 14878 13634
rect 16930 13582 16942 13634
rect 16994 13582 17006 13634
rect 23426 13582 23438 13634
rect 23490 13582 23502 13634
rect 29138 13582 29150 13634
rect 29202 13582 29214 13634
rect 38322 13582 38334 13634
rect 38386 13582 38398 13634
rect 45378 13582 45390 13634
rect 45442 13582 45454 13634
rect 7758 13570 7810 13582
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 19294 13186 19346 13198
rect 19294 13122 19346 13134
rect 19518 13186 19570 13198
rect 19518 13122 19570 13134
rect 27918 13186 27970 13198
rect 27918 13122 27970 13134
rect 28030 13186 28082 13198
rect 28030 13122 28082 13134
rect 28254 13186 28306 13198
rect 28254 13122 28306 13134
rect 28478 13186 28530 13198
rect 28478 13122 28530 13134
rect 6974 13074 7026 13086
rect 6974 13010 7026 13022
rect 19070 13074 19122 13086
rect 19070 13010 19122 13022
rect 19966 13074 20018 13086
rect 23314 13022 23326 13074
rect 23378 13022 23390 13074
rect 30706 13022 30718 13074
rect 30770 13022 30782 13074
rect 32834 13022 32846 13074
rect 32898 13022 32910 13074
rect 33394 13022 33406 13074
rect 33458 13022 33470 13074
rect 39778 13022 39790 13074
rect 39842 13022 39854 13074
rect 41906 13022 41918 13074
rect 41970 13022 41982 13074
rect 48402 13022 48414 13074
rect 48466 13022 48478 13074
rect 19966 13010 20018 13022
rect 6078 12962 6130 12974
rect 6078 12898 6130 12910
rect 7086 12962 7138 12974
rect 7086 12898 7138 12910
rect 8990 12962 9042 12974
rect 8990 12898 9042 12910
rect 9550 12962 9602 12974
rect 9550 12898 9602 12910
rect 10670 12962 10722 12974
rect 10670 12898 10722 12910
rect 11006 12962 11058 12974
rect 12798 12962 12850 12974
rect 12562 12910 12574 12962
rect 12626 12910 12638 12962
rect 11006 12898 11058 12910
rect 12798 12898 12850 12910
rect 23214 12962 23266 12974
rect 53454 12962 53506 12974
rect 23538 12910 23550 12962
rect 23602 12910 23614 12962
rect 29922 12910 29934 12962
rect 29986 12910 29998 12962
rect 36306 12910 36318 12962
rect 36370 12910 36382 12962
rect 39106 12910 39118 12962
rect 39170 12910 39182 12962
rect 45490 12910 45502 12962
rect 45554 12910 45566 12962
rect 23214 12898 23266 12910
rect 53454 12898 53506 12910
rect 53678 12962 53730 12974
rect 53678 12898 53730 12910
rect 6638 12850 6690 12862
rect 6638 12786 6690 12798
rect 9102 12850 9154 12862
rect 9102 12786 9154 12798
rect 11342 12850 11394 12862
rect 11342 12786 11394 12798
rect 11902 12850 11954 12862
rect 11902 12786 11954 12798
rect 15598 12850 15650 12862
rect 15598 12786 15650 12798
rect 18846 12850 18898 12862
rect 18846 12786 18898 12798
rect 28590 12850 28642 12862
rect 44046 12850 44098 12862
rect 54126 12850 54178 12862
rect 35522 12798 35534 12850
rect 35586 12798 35598 12850
rect 46274 12798 46286 12850
rect 46338 12798 46350 12850
rect 28590 12786 28642 12798
rect 44046 12786 44098 12798
rect 54126 12786 54178 12798
rect 5742 12738 5794 12750
rect 5742 12674 5794 12686
rect 6862 12738 6914 12750
rect 6862 12674 6914 12686
rect 7198 12738 7250 12750
rect 7198 12674 7250 12686
rect 7758 12738 7810 12750
rect 7758 12674 7810 12686
rect 9214 12738 9266 12750
rect 9214 12674 9266 12686
rect 11006 12738 11058 12750
rect 11006 12674 11058 12686
rect 14030 12738 14082 12750
rect 14030 12674 14082 12686
rect 16718 12738 16770 12750
rect 16718 12674 16770 12686
rect 17278 12738 17330 12750
rect 17278 12674 17330 12686
rect 21646 12738 21698 12750
rect 26350 12738 26402 12750
rect 23874 12686 23886 12738
rect 23938 12686 23950 12738
rect 21646 12674 21698 12686
rect 26350 12674 26402 12686
rect 36766 12738 36818 12750
rect 36766 12674 36818 12686
rect 48862 12738 48914 12750
rect 48862 12674 48914 12686
rect 53342 12738 53394 12750
rect 53342 12674 53394 12686
rect 53902 12738 53954 12750
rect 53902 12674 53954 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 23886 12402 23938 12414
rect 9762 12350 9774 12402
rect 9826 12350 9838 12402
rect 23886 12338 23938 12350
rect 33966 12402 34018 12414
rect 33966 12338 34018 12350
rect 40238 12402 40290 12414
rect 40238 12338 40290 12350
rect 54462 12402 54514 12414
rect 54462 12338 54514 12350
rect 55022 12402 55074 12414
rect 55022 12338 55074 12350
rect 10334 12290 10386 12302
rect 24334 12290 24386 12302
rect 49534 12290 49586 12302
rect 11666 12238 11678 12290
rect 11730 12238 11742 12290
rect 14354 12238 14366 12290
rect 14418 12238 14430 12290
rect 20738 12238 20750 12290
rect 20802 12238 20814 12290
rect 29922 12238 29934 12290
rect 29986 12238 29998 12290
rect 42354 12238 42366 12290
rect 42418 12238 42430 12290
rect 47618 12238 47630 12290
rect 47682 12238 47694 12290
rect 10334 12226 10386 12238
rect 24334 12226 24386 12238
rect 49534 12226 49586 12238
rect 28590 12178 28642 12190
rect 8978 12126 8990 12178
rect 9042 12126 9054 12178
rect 10994 12126 11006 12178
rect 11058 12126 11070 12178
rect 14466 12126 14478 12178
rect 14530 12126 14542 12178
rect 15250 12126 15262 12178
rect 15314 12126 15326 12178
rect 15586 12126 15598 12178
rect 15650 12126 15662 12178
rect 19954 12126 19966 12178
rect 20018 12126 20030 12178
rect 24098 12126 24110 12178
rect 24162 12126 24174 12178
rect 26674 12126 26686 12178
rect 26738 12126 26750 12178
rect 28018 12126 28030 12178
rect 28082 12126 28094 12178
rect 29138 12126 29150 12178
rect 29202 12126 29214 12178
rect 36978 12126 36990 12178
rect 37042 12126 37054 12178
rect 41570 12126 41582 12178
rect 41634 12126 41646 12178
rect 48402 12126 48414 12178
rect 48466 12126 48478 12178
rect 53666 12126 53678 12178
rect 53730 12126 53742 12178
rect 28590 12114 28642 12126
rect 23438 12066 23490 12078
rect 3938 12014 3950 12066
rect 4002 12014 4014 12066
rect 13794 12014 13806 12066
rect 13858 12014 13870 12066
rect 22866 12014 22878 12066
rect 22930 12014 22942 12066
rect 23438 12002 23490 12014
rect 26126 12066 26178 12078
rect 32050 12014 32062 12066
rect 32114 12014 32126 12066
rect 37650 12014 37662 12066
rect 37714 12014 37726 12066
rect 39778 12014 39790 12066
rect 39842 12014 39854 12066
rect 44482 12014 44494 12066
rect 44546 12014 44558 12066
rect 45490 12014 45502 12066
rect 45554 12014 45566 12066
rect 50754 12014 50766 12066
rect 50818 12014 50830 12066
rect 52882 12014 52894 12066
rect 52946 12014 52958 12066
rect 26126 12002 26178 12014
rect 10110 11954 10162 11966
rect 10110 11890 10162 11902
rect 14254 11954 14306 11966
rect 14254 11890 14306 11902
rect 24222 11954 24274 11966
rect 26686 11954 26738 11966
rect 26114 11902 26126 11954
rect 26178 11951 26190 11954
rect 26450 11951 26462 11954
rect 26178 11905 26462 11951
rect 26178 11902 26190 11905
rect 26450 11902 26462 11905
rect 26514 11902 26526 11954
rect 24222 11890 24274 11902
rect 26686 11890 26738 11902
rect 27022 11954 27074 11966
rect 27022 11890 27074 11902
rect 28366 11954 28418 11966
rect 28366 11890 28418 11902
rect 54238 11954 54290 11966
rect 54238 11890 54290 11902
rect 54574 11954 54626 11966
rect 54574 11890 54626 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 12798 11618 12850 11630
rect 12798 11554 12850 11566
rect 25006 11618 25058 11630
rect 25006 11554 25058 11566
rect 38334 11618 38386 11630
rect 38334 11554 38386 11566
rect 45726 11618 45778 11630
rect 45726 11554 45778 11566
rect 45838 11618 45890 11630
rect 45838 11554 45890 11566
rect 46062 11618 46114 11630
rect 46062 11554 46114 11566
rect 52334 11618 52386 11630
rect 52334 11554 52386 11566
rect 53566 11618 53618 11630
rect 53566 11554 53618 11566
rect 54238 11618 54290 11630
rect 54238 11554 54290 11566
rect 20414 11506 20466 11518
rect 36206 11506 36258 11518
rect 8642 11454 8654 11506
rect 8706 11454 8718 11506
rect 28354 11454 28366 11506
rect 28418 11454 28430 11506
rect 31938 11454 31950 11506
rect 32002 11454 32014 11506
rect 20414 11442 20466 11454
rect 36206 11442 36258 11454
rect 38446 11506 38498 11518
rect 38446 11442 38498 11454
rect 39118 11506 39170 11518
rect 53678 11506 53730 11518
rect 48850 11454 48862 11506
rect 48914 11454 48926 11506
rect 50978 11454 50990 11506
rect 51042 11454 51054 11506
rect 39118 11442 39170 11454
rect 53678 11442 53730 11454
rect 13022 11394 13074 11406
rect 46286 11394 46338 11406
rect 5730 11342 5742 11394
rect 5794 11342 5806 11394
rect 9986 11342 9998 11394
rect 10050 11342 10062 11394
rect 16146 11342 16158 11394
rect 16210 11342 16222 11394
rect 21970 11342 21982 11394
rect 22034 11342 22046 11394
rect 23538 11342 23550 11394
rect 23602 11342 23614 11394
rect 24210 11342 24222 11394
rect 24274 11342 24286 11394
rect 24658 11342 24670 11394
rect 24722 11342 24734 11394
rect 25554 11342 25566 11394
rect 25618 11342 25630 11394
rect 35746 11342 35758 11394
rect 35810 11342 35822 11394
rect 13022 11330 13074 11342
rect 46286 11330 46338 11342
rect 46846 11394 46898 11406
rect 46846 11330 46898 11342
rect 47518 11394 47570 11406
rect 51998 11394 52050 11406
rect 48178 11342 48190 11394
rect 48242 11342 48254 11394
rect 47518 11330 47570 11342
rect 51998 11330 52050 11342
rect 53902 11394 53954 11406
rect 53902 11330 53954 11342
rect 54126 11394 54178 11406
rect 54126 11330 54178 11342
rect 10222 11282 10274 11294
rect 22318 11282 22370 11294
rect 6514 11230 6526 11282
rect 6578 11230 6590 11282
rect 16818 11230 16830 11282
rect 16882 11230 16894 11282
rect 10222 11218 10274 11230
rect 22318 11218 22370 11230
rect 23662 11282 23714 11294
rect 46398 11282 46450 11294
rect 26226 11230 26238 11282
rect 26290 11230 26302 11282
rect 23662 11218 23714 11230
rect 46398 11218 46450 11230
rect 47406 11282 47458 11294
rect 47406 11218 47458 11230
rect 52222 11282 52274 11294
rect 52222 11218 52274 11230
rect 9214 11170 9266 11182
rect 9214 11106 9266 11118
rect 10670 11170 10722 11182
rect 10670 11106 10722 11118
rect 11902 11170 11954 11182
rect 11902 11106 11954 11118
rect 12462 11170 12514 11182
rect 12462 11106 12514 11118
rect 12686 11170 12738 11182
rect 12686 11106 12738 11118
rect 14030 11170 14082 11182
rect 14030 11106 14082 11118
rect 22206 11170 22258 11182
rect 22206 11106 22258 11118
rect 38558 11170 38610 11182
rect 38558 11106 38610 11118
rect 47182 11170 47234 11182
rect 47182 11106 47234 11118
rect 51438 11170 51490 11182
rect 51438 11106 51490 11118
rect 54910 11170 54962 11182
rect 54910 11106 54962 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 6750 10834 6802 10846
rect 6750 10770 6802 10782
rect 10110 10834 10162 10846
rect 10110 10770 10162 10782
rect 12238 10834 12290 10846
rect 12238 10770 12290 10782
rect 12798 10834 12850 10846
rect 12798 10770 12850 10782
rect 32174 10834 32226 10846
rect 32174 10770 32226 10782
rect 40014 10834 40066 10846
rect 40014 10770 40066 10782
rect 10670 10722 10722 10734
rect 10670 10658 10722 10670
rect 12126 10722 12178 10734
rect 12126 10658 12178 10670
rect 16718 10722 16770 10734
rect 16718 10658 16770 10670
rect 22878 10722 22930 10734
rect 22878 10658 22930 10670
rect 27022 10722 27074 10734
rect 27022 10658 27074 10670
rect 39454 10722 39506 10734
rect 39454 10658 39506 10670
rect 41806 10722 41858 10734
rect 41806 10658 41858 10670
rect 42814 10722 42866 10734
rect 42814 10658 42866 10670
rect 45950 10722 46002 10734
rect 45950 10658 46002 10670
rect 46622 10722 46674 10734
rect 46622 10658 46674 10670
rect 48638 10722 48690 10734
rect 56354 10670 56366 10722
rect 56418 10670 56430 10722
rect 48638 10658 48690 10670
rect 2830 10610 2882 10622
rect 2830 10546 2882 10558
rect 3166 10610 3218 10622
rect 3166 10546 3218 10558
rect 3390 10610 3442 10622
rect 3390 10546 3442 10558
rect 4398 10610 4450 10622
rect 4398 10546 4450 10558
rect 6638 10610 6690 10622
rect 6638 10546 6690 10558
rect 6974 10610 7026 10622
rect 9774 10610 9826 10622
rect 7410 10558 7422 10610
rect 7474 10558 7486 10610
rect 6974 10546 7026 10558
rect 9774 10546 9826 10558
rect 11006 10610 11058 10622
rect 32286 10610 32338 10622
rect 19058 10558 19070 10610
rect 19122 10558 19134 10610
rect 22418 10558 22430 10610
rect 22482 10558 22494 10610
rect 22642 10558 22654 10610
rect 22706 10558 22718 10610
rect 27906 10558 27918 10610
rect 27970 10558 27982 10610
rect 11006 10546 11058 10558
rect 32286 10546 32338 10558
rect 32510 10610 32562 10622
rect 32510 10546 32562 10558
rect 32734 10610 32786 10622
rect 39342 10610 39394 10622
rect 38434 10558 38446 10610
rect 38498 10558 38510 10610
rect 45154 10558 45166 10610
rect 45218 10558 45230 10610
rect 51426 10558 51438 10610
rect 51490 10558 51502 10610
rect 32734 10546 32786 10558
rect 39342 10546 39394 10558
rect 3054 10498 3106 10510
rect 3054 10434 3106 10446
rect 3950 10498 4002 10510
rect 22990 10498 23042 10510
rect 19730 10446 19742 10498
rect 19794 10446 19806 10498
rect 21858 10446 21870 10498
rect 21922 10446 21934 10498
rect 3950 10434 4002 10446
rect 22990 10434 23042 10446
rect 23326 10498 23378 10510
rect 50878 10498 50930 10510
rect 27682 10446 27694 10498
rect 27746 10446 27758 10498
rect 23326 10434 23378 10446
rect 50878 10434 50930 10446
rect 12238 10386 12290 10398
rect 7186 10334 7198 10386
rect 7250 10334 7262 10386
rect 12238 10322 12290 10334
rect 32174 10386 32226 10398
rect 32174 10322 32226 10334
rect 38446 10386 38498 10398
rect 38446 10322 38498 10334
rect 38782 10386 38834 10398
rect 38782 10322 38834 10334
rect 39454 10386 39506 10398
rect 39454 10322 39506 10334
rect 45390 10386 45442 10398
rect 45390 10322 45442 10334
rect 45614 10386 45666 10398
rect 45614 10322 45666 10334
rect 45838 10386 45890 10398
rect 45838 10322 45890 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 24446 10050 24498 10062
rect 24446 9986 24498 9998
rect 8094 9938 8146 9950
rect 19070 9938 19122 9950
rect 2594 9886 2606 9938
rect 2658 9886 2670 9938
rect 4722 9886 4734 9938
rect 4786 9886 4798 9938
rect 12226 9886 12238 9938
rect 12290 9886 12302 9938
rect 16482 9886 16494 9938
rect 16546 9886 16558 9938
rect 18610 9886 18622 9938
rect 18674 9886 18686 9938
rect 8094 9874 8146 9886
rect 19070 9874 19122 9886
rect 21982 9938 22034 9950
rect 33070 9938 33122 9950
rect 56814 9938 56866 9950
rect 32610 9886 32622 9938
rect 32674 9886 32686 9938
rect 38322 9886 38334 9938
rect 38386 9886 38398 9938
rect 40450 9886 40462 9938
rect 40514 9886 40526 9938
rect 41794 9886 41806 9938
rect 41858 9886 41870 9938
rect 43922 9886 43934 9938
rect 43986 9886 43998 9938
rect 45490 9886 45502 9938
rect 45554 9886 45566 9938
rect 47618 9886 47630 9938
rect 47682 9886 47694 9938
rect 52434 9886 52446 9938
rect 52498 9886 52510 9938
rect 53442 9886 53454 9938
rect 53506 9886 53518 9938
rect 55570 9886 55582 9938
rect 55634 9886 55646 9938
rect 21982 9874 22034 9886
rect 33070 9874 33122 9886
rect 56814 9874 56866 9886
rect 6974 9826 7026 9838
rect 1922 9774 1934 9826
rect 1986 9774 1998 9826
rect 6974 9762 7026 9774
rect 7870 9826 7922 9838
rect 7870 9762 7922 9774
rect 8542 9826 8594 9838
rect 8542 9762 8594 9774
rect 9886 9826 9938 9838
rect 9886 9762 9938 9774
rect 11006 9826 11058 9838
rect 22206 9826 22258 9838
rect 12562 9774 12574 9826
rect 12626 9774 12638 9826
rect 15698 9774 15710 9826
rect 15762 9774 15774 9826
rect 11006 9762 11058 9774
rect 22206 9762 22258 9774
rect 24670 9826 24722 9838
rect 27470 9826 27522 9838
rect 24882 9774 24894 9826
rect 24946 9774 24958 9826
rect 24670 9762 24722 9774
rect 27470 9762 27522 9774
rect 27582 9826 27634 9838
rect 27582 9762 27634 9774
rect 27806 9826 27858 9838
rect 29810 9774 29822 9826
rect 29874 9774 29886 9826
rect 37650 9774 37662 9826
rect 37714 9774 37726 9826
rect 41010 9774 41022 9826
rect 41074 9774 41086 9826
rect 48290 9774 48302 9826
rect 48354 9774 48366 9826
rect 49522 9774 49534 9826
rect 49586 9774 49598 9826
rect 56354 9774 56366 9826
rect 56418 9774 56430 9826
rect 27806 9762 27858 9774
rect 6750 9714 6802 9726
rect 6750 9650 6802 9662
rect 6862 9714 6914 9726
rect 6862 9650 6914 9662
rect 8318 9714 8370 9726
rect 8318 9650 8370 9662
rect 10782 9714 10834 9726
rect 10782 9650 10834 9662
rect 11342 9714 11394 9726
rect 11342 9650 11394 9662
rect 11902 9714 11954 9726
rect 11902 9650 11954 9662
rect 27134 9714 27186 9726
rect 30482 9662 30494 9714
rect 30546 9662 30558 9714
rect 50306 9662 50318 9714
rect 50370 9662 50382 9714
rect 27134 9650 27186 9662
rect 9326 9602 9378 9614
rect 7410 9550 7422 9602
rect 7474 9550 7486 9602
rect 9326 9538 9378 9550
rect 10222 9602 10274 9614
rect 10222 9538 10274 9550
rect 11006 9602 11058 9614
rect 24782 9602 24834 9614
rect 22530 9550 22542 9602
rect 22594 9550 22606 9602
rect 11006 9538 11058 9550
rect 24782 9538 24834 9550
rect 44382 9602 44434 9614
rect 44382 9538 44434 9550
rect 48862 9602 48914 9614
rect 48862 9538 48914 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 8206 9266 8258 9278
rect 19070 9266 19122 9278
rect 10098 9214 10110 9266
rect 10162 9214 10174 9266
rect 8206 9202 8258 9214
rect 19070 9202 19122 9214
rect 26910 9266 26962 9278
rect 26910 9202 26962 9214
rect 30718 9266 30770 9278
rect 30718 9202 30770 9214
rect 45166 9266 45218 9278
rect 45166 9202 45218 9214
rect 48078 9266 48130 9278
rect 48078 9202 48130 9214
rect 5966 9154 6018 9166
rect 8654 9154 8706 9166
rect 7634 9102 7646 9154
rect 7698 9102 7710 9154
rect 5966 9090 6018 9102
rect 8654 9090 8706 9102
rect 8878 9154 8930 9166
rect 8878 9090 8930 9102
rect 9774 9154 9826 9166
rect 48750 9154 48802 9166
rect 9986 9102 9998 9154
rect 10050 9102 10062 9154
rect 13458 9102 13470 9154
rect 13522 9102 13534 9154
rect 27458 9102 27470 9154
rect 27522 9102 27534 9154
rect 27794 9102 27806 9154
rect 27858 9102 27870 9154
rect 42578 9102 42590 9154
rect 42642 9102 42654 9154
rect 9774 9090 9826 9102
rect 48750 9090 48802 9102
rect 55358 9154 55410 9166
rect 55358 9090 55410 9102
rect 7198 9042 7250 9054
rect 4050 8990 4062 9042
rect 4114 8990 4126 9042
rect 6178 8990 6190 9042
rect 6242 8990 6254 9042
rect 7198 8978 7250 8990
rect 7422 9042 7474 9054
rect 7422 8978 7474 8990
rect 7982 9042 8034 9054
rect 16046 9042 16098 9054
rect 27134 9042 27186 9054
rect 40238 9042 40290 9054
rect 10546 8990 10558 9042
rect 10610 8990 10622 9042
rect 12786 8990 12798 9042
rect 12850 8990 12862 9042
rect 20402 8990 20414 9042
rect 20466 8990 20478 9042
rect 39442 8990 39454 9042
rect 39506 8990 39518 9042
rect 7982 8978 8034 8990
rect 16046 8978 16098 8990
rect 27134 8978 27186 8990
rect 40238 8978 40290 8990
rect 40686 9042 40738 9054
rect 41794 8990 41806 9042
rect 41858 8990 41870 9042
rect 50866 8990 50878 9042
rect 50930 8990 50942 9042
rect 40686 8978 40738 8990
rect 3278 8930 3330 8942
rect 11006 8930 11058 8942
rect 27918 8930 27970 8942
rect 3378 8878 3390 8930
rect 3442 8878 3454 8930
rect 15586 8878 15598 8930
rect 15650 8878 15662 8930
rect 23202 8878 23214 8930
rect 23266 8878 23278 8930
rect 3278 8866 3330 8878
rect 11006 8866 11058 8878
rect 27918 8866 27970 8878
rect 38670 8930 38722 8942
rect 39218 8878 39230 8930
rect 39282 8878 39294 8930
rect 44706 8878 44718 8930
rect 44770 8878 44782 8930
rect 51538 8878 51550 8930
rect 51602 8878 51614 8930
rect 38670 8866 38722 8878
rect 8990 8818 9042 8830
rect 8990 8754 9042 8766
rect 10222 8818 10274 8830
rect 10222 8754 10274 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 21758 8482 21810 8494
rect 21758 8418 21810 8430
rect 22094 8482 22146 8494
rect 22094 8418 22146 8430
rect 22878 8482 22930 8494
rect 22878 8418 22930 8430
rect 27806 8482 27858 8494
rect 27806 8418 27858 8430
rect 28030 8370 28082 8382
rect 52670 8370 52722 8382
rect 4946 8318 4958 8370
rect 5010 8318 5022 8370
rect 6514 8318 6526 8370
rect 6578 8318 6590 8370
rect 8642 8318 8654 8370
rect 8706 8318 8718 8370
rect 16594 8318 16606 8370
rect 16658 8318 16670 8370
rect 18722 8318 18734 8370
rect 18786 8318 18798 8370
rect 24770 8318 24782 8370
rect 24834 8318 24846 8370
rect 26898 8318 26910 8370
rect 26962 8318 26974 8370
rect 51874 8318 51886 8370
rect 51938 8318 51950 8370
rect 28030 8306 28082 8318
rect 52670 8306 52722 8318
rect 9662 8258 9714 8270
rect 2146 8206 2158 8258
rect 2210 8206 2222 8258
rect 5730 8206 5742 8258
rect 5794 8206 5806 8258
rect 9662 8194 9714 8206
rect 10222 8258 10274 8270
rect 10222 8194 10274 8206
rect 11006 8258 11058 8270
rect 11566 8258 11618 8270
rect 11330 8206 11342 8258
rect 11394 8206 11406 8258
rect 11006 8194 11058 8206
rect 11566 8194 11618 8206
rect 11790 8258 11842 8270
rect 20862 8258 20914 8270
rect 15810 8206 15822 8258
rect 15874 8206 15886 8258
rect 11790 8194 11842 8206
rect 20862 8194 20914 8206
rect 21870 8258 21922 8270
rect 53566 8258 53618 8270
rect 22306 8206 22318 8258
rect 22370 8206 22382 8258
rect 23986 8206 23998 8258
rect 24050 8206 24062 8258
rect 44594 8206 44606 8258
rect 44658 8206 44670 8258
rect 48962 8206 48974 8258
rect 49026 8206 49038 8258
rect 49746 8206 49758 8258
rect 49810 8206 49822 8258
rect 21870 8194 21922 8206
rect 53566 8194 53618 8206
rect 53790 8258 53842 8270
rect 53790 8194 53842 8206
rect 54014 8258 54066 8270
rect 54014 8194 54066 8206
rect 54126 8258 54178 8270
rect 54126 8194 54178 8206
rect 10110 8146 10162 8158
rect 2818 8094 2830 8146
rect 2882 8094 2894 8146
rect 10110 8082 10162 8094
rect 12014 8146 12066 8158
rect 42466 8094 42478 8146
rect 42530 8094 42542 8146
rect 12014 8082 12066 8094
rect 9214 8034 9266 8046
rect 9214 7970 9266 7982
rect 9886 8034 9938 8046
rect 9886 7970 9938 7982
rect 12126 8034 12178 8046
rect 12126 7970 12178 7982
rect 19182 8034 19234 8046
rect 19182 7970 19234 7982
rect 20638 8034 20690 8046
rect 20638 7970 20690 7982
rect 20750 8034 20802 8046
rect 20750 7970 20802 7982
rect 22990 8034 23042 8046
rect 22990 7970 23042 7982
rect 23102 8034 23154 8046
rect 38782 8034 38834 8046
rect 27458 7982 27470 8034
rect 27522 7982 27534 8034
rect 23102 7970 23154 7982
rect 38782 7970 38834 7982
rect 45502 8034 45554 8046
rect 45502 7970 45554 7982
rect 47182 8034 47234 8046
rect 47182 7970 47234 7982
rect 54126 8034 54178 8046
rect 54126 7970 54178 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 2830 7698 2882 7710
rect 2830 7634 2882 7646
rect 15934 7698 15986 7710
rect 15934 7634 15986 7646
rect 30494 7698 30546 7710
rect 30494 7634 30546 7646
rect 51774 7698 51826 7710
rect 51774 7634 51826 7646
rect 55694 7698 55746 7710
rect 55694 7634 55746 7646
rect 3166 7586 3218 7598
rect 22766 7586 22818 7598
rect 3938 7534 3950 7586
rect 4002 7534 4014 7586
rect 14690 7534 14702 7586
rect 14754 7534 14766 7586
rect 3166 7522 3218 7534
rect 22766 7522 22818 7534
rect 22990 7586 23042 7598
rect 22990 7522 23042 7534
rect 24670 7586 24722 7598
rect 24670 7522 24722 7534
rect 26238 7586 26290 7598
rect 50430 7586 50482 7598
rect 43250 7534 43262 7586
rect 43314 7534 43326 7586
rect 54450 7534 54462 7586
rect 54514 7534 54526 7586
rect 26238 7522 26290 7534
rect 50430 7522 50482 7534
rect 2606 7474 2658 7486
rect 2606 7410 2658 7422
rect 2830 7474 2882 7486
rect 8978 7422 8990 7474
rect 9042 7422 9054 7474
rect 10882 7422 10894 7474
rect 10946 7422 10958 7474
rect 15474 7422 15486 7474
rect 15538 7422 15550 7474
rect 19170 7422 19182 7474
rect 19234 7422 19246 7474
rect 26562 7422 26574 7474
rect 26626 7422 26638 7474
rect 29922 7422 29934 7474
rect 29986 7422 29998 7474
rect 38210 7422 38222 7474
rect 38274 7422 38286 7474
rect 39330 7422 39342 7474
rect 39394 7422 39406 7474
rect 39778 7422 39790 7474
rect 39842 7422 39854 7474
rect 42466 7422 42478 7474
rect 42530 7422 42542 7474
rect 55234 7422 55246 7474
rect 55298 7422 55310 7474
rect 2830 7410 2882 7422
rect 23662 7362 23714 7374
rect 10770 7310 10782 7362
rect 10834 7310 10846 7362
rect 12562 7310 12574 7362
rect 12626 7310 12638 7362
rect 19954 7310 19966 7362
rect 20018 7310 20030 7362
rect 22082 7310 22094 7362
rect 22146 7310 22158 7362
rect 22642 7310 22654 7362
rect 22706 7310 22718 7362
rect 23662 7298 23714 7310
rect 24558 7362 24610 7374
rect 24558 7298 24610 7310
rect 25566 7362 25618 7374
rect 38558 7362 38610 7374
rect 27122 7310 27134 7362
rect 27186 7310 27198 7362
rect 29250 7310 29262 7362
rect 29314 7310 29326 7362
rect 38322 7310 38334 7362
rect 38386 7310 38398 7362
rect 25566 7298 25618 7310
rect 38558 7298 38610 7310
rect 39118 7362 39170 7374
rect 39118 7298 39170 7310
rect 41918 7362 41970 7374
rect 45378 7310 45390 7362
rect 45442 7310 45454 7362
rect 52322 7310 52334 7362
rect 52386 7310 52398 7362
rect 41918 7298 41970 7310
rect 24446 7250 24498 7262
rect 10210 7198 10222 7250
rect 10274 7198 10286 7250
rect 24446 7186 24498 7198
rect 26574 7250 26626 7262
rect 26574 7186 26626 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 27694 6914 27746 6926
rect 11890 6862 11902 6914
rect 11954 6862 11966 6914
rect 27694 6850 27746 6862
rect 12238 6802 12290 6814
rect 9202 6750 9214 6802
rect 9266 6750 9278 6802
rect 11330 6750 11342 6802
rect 11394 6750 11406 6802
rect 12238 6738 12290 6750
rect 22654 6802 22706 6814
rect 26798 6802 26850 6814
rect 53342 6802 53394 6814
rect 23874 6750 23886 6802
rect 23938 6750 23950 6802
rect 26002 6750 26014 6802
rect 26066 6750 26078 6802
rect 38322 6750 38334 6802
rect 38386 6750 38398 6802
rect 40450 6750 40462 6802
rect 40514 6750 40526 6802
rect 49074 6750 49086 6802
rect 49138 6750 49150 6802
rect 50418 6750 50430 6802
rect 50482 6750 50494 6802
rect 52546 6750 52558 6802
rect 52610 6750 52622 6802
rect 22654 6738 22706 6750
rect 26798 6738 26850 6750
rect 53342 6738 53394 6750
rect 2270 6690 2322 6702
rect 2270 6626 2322 6638
rect 2718 6690 2770 6702
rect 2718 6626 2770 6638
rect 4174 6690 4226 6702
rect 12462 6690 12514 6702
rect 27470 6690 27522 6702
rect 8530 6638 8542 6690
rect 8594 6638 8606 6690
rect 23202 6638 23214 6690
rect 23266 6638 23278 6690
rect 27234 6638 27246 6690
rect 27298 6638 27310 6690
rect 4174 6626 4226 6638
rect 12462 6626 12514 6638
rect 27470 6626 27522 6638
rect 27806 6690 27858 6702
rect 37650 6638 37662 6690
rect 37714 6638 37726 6690
rect 46274 6638 46286 6690
rect 46338 6638 46350 6690
rect 46946 6638 46958 6690
rect 47010 6638 47022 6690
rect 49634 6638 49646 6690
rect 49698 6638 49710 6690
rect 27806 6626 27858 6638
rect 3726 6578 3778 6590
rect 3726 6514 3778 6526
rect 2830 6466 2882 6478
rect 2830 6402 2882 6414
rect 22094 6466 22146 6478
rect 22094 6402 22146 6414
rect 40910 6466 40962 6478
rect 40910 6402 40962 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 11790 6130 11842 6142
rect 11790 6066 11842 6078
rect 22430 6130 22482 6142
rect 22430 6066 22482 6078
rect 26238 6130 26290 6142
rect 26238 6066 26290 6078
rect 40014 6130 40066 6142
rect 40014 6066 40066 6078
rect 49422 6130 49474 6142
rect 49422 6066 49474 6078
rect 52782 6130 52834 6142
rect 52782 6066 52834 6078
rect 11902 6018 11954 6030
rect 3938 5966 3950 6018
rect 4002 5966 4014 6018
rect 11902 5954 11954 5966
rect 12126 6018 12178 6030
rect 39230 6018 39282 6030
rect 19842 5966 19854 6018
rect 19906 5966 19918 6018
rect 12126 5954 12178 5966
rect 39230 5954 39282 5966
rect 39790 6018 39842 6030
rect 54114 5966 54126 6018
rect 54178 5966 54190 6018
rect 39790 5954 39842 5966
rect 11454 5906 11506 5918
rect 4722 5854 4734 5906
rect 4786 5854 4798 5906
rect 19170 5854 19182 5906
rect 19234 5854 19246 5906
rect 53330 5854 53342 5906
rect 53394 5854 53406 5906
rect 11454 5842 11506 5854
rect 1810 5742 1822 5794
rect 1874 5742 1886 5794
rect 21970 5742 21982 5794
rect 22034 5742 22046 5794
rect 56242 5742 56254 5794
rect 56306 5742 56318 5794
rect 40126 5682 40178 5694
rect 40126 5618 40178 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 41234 5182 41246 5234
rect 41298 5182 41310 5234
rect 43362 5182 43374 5234
rect 43426 5182 43438 5234
rect 55346 5182 55358 5234
rect 55410 5182 55422 5234
rect 43934 5122 43986 5134
rect 40562 5070 40574 5122
rect 40626 5070 40638 5122
rect 56130 5070 56142 5122
rect 56194 5070 56206 5122
rect 43934 5058 43986 5070
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 2482 3614 2494 3666
rect 2546 3614 2558 3666
rect 22418 3614 22430 3666
rect 22482 3614 22494 3666
rect 45602 3614 45614 3666
rect 45666 3614 45678 3666
rect 1810 3502 1822 3554
rect 1874 3502 1886 3554
rect 21970 3502 21982 3554
rect 22034 3502 22046 3554
rect 44930 3502 44942 3554
rect 44994 3502 45006 3554
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 5406 56590 5458 56642
rect 6414 56590 6466 56642
rect 26910 56590 26962 56642
rect 27806 56590 27858 56642
rect 49086 56590 49138 56642
rect 49982 56590 50034 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 5070 56030 5122 56082
rect 5742 56030 5794 56082
rect 27246 56030 27298 56082
rect 49310 56030 49362 56082
rect 6414 55918 6466 55970
rect 27806 55918 27858 55970
rect 49982 55918 50034 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 8318 52110 8370 52162
rect 9102 52110 9154 52162
rect 8430 51886 8482 51938
rect 8542 51886 8594 51938
rect 19518 51886 19570 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 19294 51438 19346 51490
rect 41582 51438 41634 51490
rect 8990 51326 9042 51378
rect 9774 51326 9826 51378
rect 18510 51326 18562 51378
rect 33966 51326 34018 51378
rect 45950 51326 46002 51378
rect 49534 51326 49586 51378
rect 4958 51214 5010 51266
rect 13246 51214 13298 51266
rect 21422 51214 21474 51266
rect 21982 51214 22034 51266
rect 26238 51214 26290 51266
rect 34750 51214 34802 51266
rect 36878 51214 36930 51266
rect 37438 51214 37490 51266
rect 46622 51214 46674 51266
rect 48750 51214 48802 51266
rect 50318 51214 50370 51266
rect 52446 51214 52498 51266
rect 53006 51214 53058 51266
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 2046 50654 2098 50706
rect 4174 50654 4226 50706
rect 9438 50654 9490 50706
rect 12910 50654 12962 50706
rect 13694 50654 13746 50706
rect 27246 50654 27298 50706
rect 40798 50654 40850 50706
rect 42926 50654 42978 50706
rect 4958 50542 5010 50594
rect 6526 50542 6578 50594
rect 10110 50542 10162 50594
rect 16606 50542 16658 50594
rect 24446 50542 24498 50594
rect 40014 50542 40066 50594
rect 7310 50430 7362 50482
rect 10782 50430 10834 50482
rect 15822 50430 15874 50482
rect 17054 50430 17106 50482
rect 25118 50430 25170 50482
rect 34862 50430 34914 50482
rect 39454 50430 39506 50482
rect 50318 50430 50370 50482
rect 54238 50430 54290 50482
rect 21646 50318 21698 50370
rect 27694 50318 27746 50370
rect 37662 50318 37714 50370
rect 48974 50318 49026 50370
rect 53342 50318 53394 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 8654 49982 8706 50034
rect 9886 49982 9938 50034
rect 11678 49982 11730 50034
rect 23326 49982 23378 50034
rect 42702 49982 42754 50034
rect 47630 49982 47682 50034
rect 9774 49870 9826 49922
rect 12462 49870 12514 49922
rect 12686 49870 12738 49922
rect 13918 49870 13970 49922
rect 16382 49870 16434 49922
rect 20750 49870 20802 49922
rect 25790 49870 25842 49922
rect 41694 49870 41746 49922
rect 47742 49870 47794 49922
rect 4286 49758 4338 49810
rect 8318 49758 8370 49810
rect 8654 49758 8706 49810
rect 8990 49758 9042 49810
rect 10110 49758 10162 49810
rect 11902 49758 11954 49810
rect 13358 49758 13410 49810
rect 19966 49758 20018 49810
rect 27694 49758 27746 49810
rect 36878 49758 36930 49810
rect 42254 49758 42306 49810
rect 42814 49758 42866 49810
rect 43262 49758 43314 49810
rect 43486 49758 43538 49810
rect 46958 49758 47010 49810
rect 51102 49758 51154 49810
rect 56142 49758 56194 49810
rect 4958 49646 5010 49698
rect 7086 49646 7138 49698
rect 12798 49646 12850 49698
rect 22878 49646 22930 49698
rect 24894 49646 24946 49698
rect 25678 49646 25730 49698
rect 26462 49646 26514 49698
rect 27134 49646 27186 49698
rect 28366 49646 28418 49698
rect 30494 49646 30546 49698
rect 30942 49646 30994 49698
rect 37886 49646 37938 49698
rect 44046 49646 44098 49698
rect 46174 49646 46226 49698
rect 51886 49646 51938 49698
rect 54014 49646 54066 49698
rect 55358 49646 55410 49698
rect 11566 49534 11618 49586
rect 13582 49534 13634 49586
rect 13806 49534 13858 49586
rect 24782 49534 24834 49586
rect 26014 49534 26066 49586
rect 42926 49534 42978 49586
rect 47518 49534 47570 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 12574 49198 12626 49250
rect 22094 49198 22146 49250
rect 22318 49198 22370 49250
rect 28366 49198 28418 49250
rect 45838 49198 45890 49250
rect 15150 49086 15202 49138
rect 17278 49086 17330 49138
rect 20750 49086 20802 49138
rect 21870 49086 21922 49138
rect 22990 49086 23042 49138
rect 36318 49086 36370 49138
rect 36766 49086 36818 49138
rect 37550 49086 37602 49138
rect 39678 49086 39730 49138
rect 41806 49086 41858 49138
rect 43934 49086 43986 49138
rect 52446 49086 52498 49138
rect 56478 49086 56530 49138
rect 7310 48974 7362 49026
rect 7534 48974 7586 49026
rect 12350 48974 12402 49026
rect 14366 48974 14418 49026
rect 17950 48974 18002 49026
rect 21646 48974 21698 49026
rect 25902 48974 25954 49026
rect 26350 48974 26402 49026
rect 26686 48974 26738 49026
rect 30270 48974 30322 49026
rect 30942 48974 30994 49026
rect 40350 48974 40402 49026
rect 41022 48974 41074 49026
rect 45838 48974 45890 49026
rect 49534 48974 49586 49026
rect 53566 48974 53618 49026
rect 8766 48862 8818 48914
rect 18622 48862 18674 48914
rect 25118 48862 25170 48914
rect 26574 48862 26626 48914
rect 27022 48862 27074 48914
rect 28702 48862 28754 48914
rect 30046 48862 30098 48914
rect 45502 48862 45554 48914
rect 48974 48862 49026 48914
rect 50318 48862 50370 48914
rect 54350 48862 54402 48914
rect 56926 48862 56978 48914
rect 7870 48750 7922 48802
rect 8542 48750 8594 48802
rect 8654 48750 8706 48802
rect 12910 48750 12962 48802
rect 22206 48750 22258 48802
rect 27806 48750 27858 48802
rect 28478 48750 28530 48802
rect 33854 48750 33906 48802
rect 35198 48750 35250 48802
rect 47182 48750 47234 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 18734 48414 18786 48466
rect 20974 48414 21026 48466
rect 24670 48414 24722 48466
rect 36990 48414 37042 48466
rect 41470 48414 41522 48466
rect 7310 48302 7362 48354
rect 8542 48302 8594 48354
rect 24446 48302 24498 48354
rect 32510 48302 32562 48354
rect 34414 48302 34466 48354
rect 44718 48302 44770 48354
rect 48078 48302 48130 48354
rect 7422 48190 7474 48242
rect 7646 48190 7698 48242
rect 9662 48190 9714 48242
rect 12574 48190 12626 48242
rect 12798 48190 12850 48242
rect 13134 48190 13186 48242
rect 13918 48190 13970 48242
rect 24334 48190 24386 48242
rect 27358 48190 27410 48242
rect 32734 48190 32786 48242
rect 33742 48190 33794 48242
rect 37886 48190 37938 48242
rect 44046 48190 44098 48242
rect 48750 48190 48802 48242
rect 49534 48190 49586 48242
rect 8542 48078 8594 48130
rect 12910 48078 12962 48130
rect 14030 48078 14082 48130
rect 17614 48078 17666 48130
rect 25678 48078 25730 48130
rect 31726 48078 31778 48130
rect 36542 48078 36594 48130
rect 38670 48078 38722 48130
rect 40798 48078 40850 48130
rect 44494 48078 44546 48130
rect 51550 48078 51602 48130
rect 7758 47966 7810 48018
rect 8766 47966 8818 48018
rect 14254 47966 14306 48018
rect 25790 47966 25842 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 21646 47630 21698 47682
rect 37774 47630 37826 47682
rect 38222 47630 38274 47682
rect 7870 47518 7922 47570
rect 22206 47518 22258 47570
rect 24334 47518 24386 47570
rect 27918 47518 27970 47570
rect 28814 47518 28866 47570
rect 34638 47518 34690 47570
rect 36766 47518 36818 47570
rect 37998 47518 38050 47570
rect 45502 47518 45554 47570
rect 47966 47518 48018 47570
rect 50094 47518 50146 47570
rect 7646 47406 7698 47458
rect 8654 47406 8706 47458
rect 8878 47406 8930 47458
rect 9102 47406 9154 47458
rect 12238 47406 12290 47458
rect 12686 47406 12738 47458
rect 12798 47406 12850 47458
rect 14142 47406 14194 47458
rect 21982 47406 22034 47458
rect 23214 47406 23266 47458
rect 24222 47406 24274 47458
rect 25118 47406 25170 47458
rect 30718 47406 30770 47458
rect 31054 47406 31106 47458
rect 31614 47406 31666 47458
rect 32174 47406 32226 47458
rect 33854 47406 33906 47458
rect 37550 47406 37602 47458
rect 47182 47406 47234 47458
rect 54014 47406 54066 47458
rect 55134 47406 55186 47458
rect 8430 47294 8482 47346
rect 10110 47294 10162 47346
rect 10446 47294 10498 47346
rect 12462 47294 12514 47346
rect 16830 47294 16882 47346
rect 23438 47294 23490 47346
rect 24110 47294 24162 47346
rect 25790 47294 25842 47346
rect 28478 47294 28530 47346
rect 28702 47294 28754 47346
rect 29486 47294 29538 47346
rect 30830 47294 30882 47346
rect 31838 47294 31890 47346
rect 38334 47294 38386 47346
rect 39118 47294 39170 47346
rect 45614 47294 45666 47346
rect 45838 47294 45890 47346
rect 52110 47294 52162 47346
rect 53454 47294 53506 47346
rect 55022 47294 55074 47346
rect 7310 47182 7362 47234
rect 9214 47182 9266 47234
rect 11902 47182 11954 47234
rect 19518 47182 19570 47234
rect 20750 47182 20802 47234
rect 30270 47182 30322 47234
rect 31950 47182 32002 47234
rect 50542 47182 50594 47234
rect 52670 47182 52722 47234
rect 54014 47182 54066 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 17614 46846 17666 46898
rect 37102 46846 37154 46898
rect 47182 46846 47234 46898
rect 54574 46846 54626 46898
rect 3502 46734 3554 46786
rect 5742 46734 5794 46786
rect 8990 46734 9042 46786
rect 16942 46734 16994 46786
rect 24670 46734 24722 46786
rect 25678 46734 25730 46786
rect 27806 46734 27858 46786
rect 29150 46734 29202 46786
rect 38334 46734 38386 46786
rect 41694 46734 41746 46786
rect 42030 46734 42082 46786
rect 45166 46734 45218 46786
rect 48526 46734 48578 46786
rect 5070 46622 5122 46674
rect 8542 46622 8594 46674
rect 8654 46622 8706 46674
rect 8878 46622 8930 46674
rect 9886 46622 9938 46674
rect 16158 46622 16210 46674
rect 18398 46622 18450 46674
rect 26014 46622 26066 46674
rect 27470 46622 27522 46674
rect 28478 46622 28530 46674
rect 41582 46622 41634 46674
rect 42366 46622 42418 46674
rect 45838 46622 45890 46674
rect 46398 46622 46450 46674
rect 47070 46622 47122 46674
rect 47742 46622 47794 46674
rect 48414 46622 48466 46674
rect 51214 46622 51266 46674
rect 7870 46510 7922 46562
rect 10558 46510 10610 46562
rect 12686 46510 12738 46562
rect 13246 46510 13298 46562
rect 15374 46510 15426 46562
rect 22878 46510 22930 46562
rect 24782 46510 24834 46562
rect 25790 46510 25842 46562
rect 26126 46510 26178 46562
rect 26910 46510 26962 46562
rect 31278 46510 31330 46562
rect 31726 46510 31778 46562
rect 40798 46510 40850 46562
rect 43038 46510 43090 46562
rect 49534 46510 49586 46562
rect 51998 46510 52050 46562
rect 54126 46510 54178 46562
rect 24894 46398 24946 46450
rect 42590 46398 42642 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 10334 46062 10386 46114
rect 10782 46062 10834 46114
rect 21758 46062 21810 46114
rect 25902 46062 25954 46114
rect 29822 46062 29874 46114
rect 30158 46062 30210 46114
rect 2830 45950 2882 46002
rect 4958 45950 5010 46002
rect 9214 45950 9266 46002
rect 12910 45950 12962 46002
rect 13582 45950 13634 46002
rect 17390 45950 17442 46002
rect 18734 45950 18786 46002
rect 20862 45950 20914 46002
rect 21870 45950 21922 46002
rect 22878 45950 22930 46002
rect 30830 45950 30882 46002
rect 38334 45950 38386 46002
rect 40462 45950 40514 46002
rect 43934 45950 43986 46002
rect 48414 45950 48466 46002
rect 48974 45950 49026 46002
rect 2046 45838 2098 45890
rect 10446 45838 10498 45890
rect 10670 45838 10722 45890
rect 14478 45838 14530 45890
rect 18062 45838 18114 45890
rect 22094 45838 22146 45890
rect 22318 45838 22370 45890
rect 25566 45838 25618 45890
rect 26126 45838 26178 45890
rect 26798 45838 26850 45890
rect 29934 45838 29986 45890
rect 33630 45838 33682 45890
rect 37662 45838 37714 45890
rect 41022 45838 41074 45890
rect 45614 45838 45666 45890
rect 15262 45726 15314 45778
rect 25790 45726 25842 45778
rect 32958 45726 33010 45778
rect 41806 45726 41858 45778
rect 46286 45726 46338 45778
rect 52110 45726 52162 45778
rect 5630 45614 5682 45666
rect 8094 45614 8146 45666
rect 22206 45614 22258 45666
rect 28142 45614 28194 45666
rect 28814 45614 28866 45666
rect 29822 45614 29874 45666
rect 34190 45614 34242 45666
rect 44382 45614 44434 45666
rect 49758 45614 49810 45666
rect 54014 45614 54066 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 4958 45278 5010 45330
rect 10558 45278 10610 45330
rect 13806 45278 13858 45330
rect 16382 45278 16434 45330
rect 17726 45278 17778 45330
rect 23214 45278 23266 45330
rect 26686 45278 26738 45330
rect 40798 45278 40850 45330
rect 2718 45166 2770 45218
rect 7310 45166 7362 45218
rect 9774 45166 9826 45218
rect 14030 45166 14082 45218
rect 20638 45166 20690 45218
rect 28366 45166 28418 45218
rect 30942 45166 30994 45218
rect 42366 45166 42418 45218
rect 50318 45166 50370 45218
rect 53790 45166 53842 45218
rect 9998 45054 10050 45106
rect 10222 45054 10274 45106
rect 10446 45054 10498 45106
rect 19966 45054 20018 45106
rect 25790 45054 25842 45106
rect 26014 45054 26066 45106
rect 26238 45054 26290 45106
rect 28142 45054 28194 45106
rect 30270 45054 30322 45106
rect 30606 45054 30658 45106
rect 31054 45054 31106 45106
rect 31278 45054 31330 45106
rect 35310 45054 35362 45106
rect 41582 45054 41634 45106
rect 42030 45054 42082 45106
rect 43822 45054 43874 45106
rect 49646 45054 49698 45106
rect 53006 45054 53058 45106
rect 13694 44942 13746 44994
rect 22766 44942 22818 44994
rect 26126 44942 26178 44994
rect 35982 44942 36034 44994
rect 38110 44942 38162 44994
rect 38558 44942 38610 44994
rect 41806 44942 41858 44994
rect 42254 44942 42306 44994
rect 44494 44942 44546 44994
rect 46622 44942 46674 44994
rect 47070 44942 47122 44994
rect 52446 44942 52498 44994
rect 55918 44942 55970 44994
rect 56366 44942 56418 44994
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 9774 44494 9826 44546
rect 25454 44494 25506 44546
rect 26910 44494 26962 44546
rect 27134 44494 27186 44546
rect 27246 44494 27298 44546
rect 29710 44494 29762 44546
rect 30718 44494 30770 44546
rect 2606 44382 2658 44434
rect 4734 44382 4786 44434
rect 5854 44382 5906 44434
rect 7198 44382 7250 44434
rect 9326 44382 9378 44434
rect 16606 44382 16658 44434
rect 17166 44382 17218 44434
rect 24670 44382 24722 44434
rect 28926 44382 28978 44434
rect 29934 44382 29986 44434
rect 48526 44382 48578 44434
rect 50878 44382 50930 44434
rect 52670 44382 52722 44434
rect 54686 44382 54738 44434
rect 1934 44270 1986 44322
rect 6414 44270 6466 44322
rect 10110 44270 10162 44322
rect 10334 44270 10386 44322
rect 13806 44270 13858 44322
rect 20862 44270 20914 44322
rect 21758 44270 21810 44322
rect 25902 44270 25954 44322
rect 26014 44270 26066 44322
rect 26238 44270 26290 44322
rect 30158 44270 30210 44322
rect 30830 44270 30882 44322
rect 31054 44270 31106 44322
rect 48078 44270 48130 44322
rect 49086 44270 49138 44322
rect 54014 44270 54066 44322
rect 54462 44270 54514 44322
rect 9886 44158 9938 44210
rect 14478 44158 14530 44210
rect 22542 44158 22594 44210
rect 26798 44158 26850 44210
rect 29598 44158 29650 44210
rect 36206 44158 36258 44210
rect 44606 44158 44658 44210
rect 46398 44158 46450 44210
rect 47406 44158 47458 44210
rect 48974 44158 49026 44210
rect 53454 44158 53506 44210
rect 55134 44158 55186 44210
rect 19294 44046 19346 44098
rect 33966 44046 34018 44098
rect 42366 44046 42418 44098
rect 45838 44046 45890 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 9886 43710 9938 43762
rect 13806 43710 13858 43762
rect 31166 43710 31218 43762
rect 48414 43710 48466 43762
rect 2830 43598 2882 43650
rect 5854 43598 5906 43650
rect 19070 43598 19122 43650
rect 21646 43598 21698 43650
rect 28590 43598 28642 43650
rect 39678 43598 39730 43650
rect 46958 43598 47010 43650
rect 50654 43598 50706 43650
rect 56254 43598 56306 43650
rect 8318 43486 8370 43538
rect 10222 43486 10274 43538
rect 15262 43486 15314 43538
rect 15710 43486 15762 43538
rect 18398 43486 18450 43538
rect 25902 43486 25954 43538
rect 26126 43486 26178 43538
rect 27918 43486 27970 43538
rect 35086 43486 35138 43538
rect 42142 43486 42194 43538
rect 51214 43486 51266 43538
rect 10782 43374 10834 43426
rect 21198 43374 21250 43426
rect 30718 43374 30770 43426
rect 35758 43374 35810 43426
rect 40238 43374 40290 43426
rect 49422 43374 49474 43426
rect 9886 43262 9938 43314
rect 9998 43262 10050 43314
rect 15486 43262 15538 43314
rect 15934 43262 15986 43314
rect 16046 43262 16098 43314
rect 26014 43262 26066 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 9102 42926 9154 42978
rect 9774 42926 9826 42978
rect 14254 42926 14306 42978
rect 14590 42926 14642 42978
rect 2830 42814 2882 42866
rect 4958 42814 5010 42866
rect 8878 42814 8930 42866
rect 12910 42814 12962 42866
rect 15374 42814 15426 42866
rect 18846 42814 18898 42866
rect 23550 42814 23602 42866
rect 34414 42814 34466 42866
rect 36542 42814 36594 42866
rect 39454 42814 39506 42866
rect 41582 42814 41634 42866
rect 42366 42814 42418 42866
rect 46286 42814 46338 42866
rect 48414 42814 48466 42866
rect 48974 42814 49026 42866
rect 51102 42814 51154 42866
rect 52334 42814 52386 42866
rect 2158 42702 2210 42754
rect 6078 42702 6130 42754
rect 9998 42702 10050 42754
rect 14814 42702 14866 42754
rect 18286 42702 18338 42754
rect 26462 42702 26514 42754
rect 33630 42702 33682 42754
rect 38782 42702 38834 42754
rect 42254 42702 42306 42754
rect 42590 42702 42642 42754
rect 42814 42702 42866 42754
rect 44718 42702 44770 42754
rect 45614 42702 45666 42754
rect 51886 42702 51938 42754
rect 6750 42590 6802 42642
rect 10782 42590 10834 42642
rect 17502 42590 17554 42642
rect 25678 42590 25730 42642
rect 9326 42478 9378 42530
rect 13582 42478 13634 42530
rect 20302 42478 20354 42530
rect 20862 42478 20914 42530
rect 37550 42478 37602 42530
rect 38110 42478 38162 42530
rect 42702 42478 42754 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 6862 42142 6914 42194
rect 16494 42142 16546 42194
rect 25790 42142 25842 42194
rect 26574 42142 26626 42194
rect 44942 42142 44994 42194
rect 53342 42142 53394 42194
rect 2718 42030 2770 42082
rect 20190 42030 20242 42082
rect 26014 42030 26066 42082
rect 32622 42030 32674 42082
rect 34302 42030 34354 42082
rect 34750 42030 34802 42082
rect 37214 42030 37266 42082
rect 4398 41918 4450 41970
rect 5182 41918 5234 41970
rect 5406 41918 5458 41970
rect 15038 41918 15090 41970
rect 15822 41918 15874 41970
rect 19406 41918 19458 41970
rect 29262 41918 29314 41970
rect 36542 41918 36594 41970
rect 41582 41918 41634 41970
rect 42366 41918 42418 41970
rect 50094 41918 50146 41970
rect 50766 41918 50818 41970
rect 4958 41806 5010 41858
rect 5630 41806 5682 41858
rect 10334 41806 10386 41858
rect 22318 41806 22370 41858
rect 22766 41806 22818 41858
rect 25678 41806 25730 41858
rect 29934 41806 29986 41858
rect 32062 41806 32114 41858
rect 39342 41806 39394 41858
rect 44494 41806 44546 41858
rect 52894 41806 52946 41858
rect 6078 41694 6130 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 22094 41358 22146 41410
rect 23774 41358 23826 41410
rect 35198 41358 35250 41410
rect 35534 41358 35586 41410
rect 2606 41246 2658 41298
rect 4734 41246 4786 41298
rect 5742 41246 5794 41298
rect 11230 41246 11282 41298
rect 20638 41246 20690 41298
rect 21870 41246 21922 41298
rect 32286 41246 32338 41298
rect 34414 41246 34466 41298
rect 35310 41246 35362 41298
rect 1934 41134 1986 41186
rect 8430 41134 8482 41186
rect 12350 41134 12402 41186
rect 17726 41134 17778 41186
rect 21646 41134 21698 41186
rect 22318 41134 22370 41186
rect 22990 41134 23042 41186
rect 31614 41134 31666 41186
rect 35758 41134 35810 41186
rect 42478 41134 42530 41186
rect 9102 41022 9154 41074
rect 11790 41022 11842 41074
rect 18510 41022 18562 41074
rect 22430 41022 22482 41074
rect 22654 41022 22706 41074
rect 22878 41022 22930 41074
rect 23214 41022 23266 41074
rect 23326 41022 23378 41074
rect 30158 41022 30210 41074
rect 40910 41022 40962 41074
rect 13694 40910 13746 40962
rect 24334 40910 24386 40962
rect 27022 40910 27074 40962
rect 35646 40910 35698 40962
rect 38110 40910 38162 40962
rect 44382 40910 44434 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 9774 40574 9826 40626
rect 11678 40574 11730 40626
rect 18062 40574 18114 40626
rect 36990 40574 37042 40626
rect 54126 40574 54178 40626
rect 5854 40462 5906 40514
rect 13022 40462 13074 40514
rect 29262 40462 29314 40514
rect 34414 40462 34466 40514
rect 38558 40462 38610 40514
rect 12350 40350 12402 40402
rect 19070 40350 19122 40402
rect 21086 40350 21138 40402
rect 25678 40350 25730 40402
rect 26686 40350 26738 40402
rect 27246 40350 27298 40402
rect 33630 40350 33682 40402
rect 37886 40350 37938 40402
rect 46622 40350 46674 40402
rect 49534 40350 49586 40402
rect 50878 40350 50930 40402
rect 8094 40238 8146 40290
rect 15150 40238 15202 40290
rect 23550 40238 23602 40290
rect 36542 40238 36594 40290
rect 40686 40238 40738 40290
rect 43710 40238 43762 40290
rect 45838 40238 45890 40290
rect 51550 40238 51602 40290
rect 53678 40238 53730 40290
rect 49758 40126 49810 40178
rect 50094 40126 50146 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 10446 39678 10498 39730
rect 12462 39678 12514 39730
rect 19966 39678 20018 39730
rect 22990 39678 23042 39730
rect 25118 39678 25170 39730
rect 25678 39678 25730 39730
rect 27806 39678 27858 39730
rect 32510 39678 32562 39730
rect 43822 39678 43874 39730
rect 47630 39678 47682 39730
rect 53678 39678 53730 39730
rect 7646 39566 7698 39618
rect 17166 39566 17218 39618
rect 22318 39566 22370 39618
rect 28590 39566 28642 39618
rect 29710 39566 29762 39618
rect 32958 39566 33010 39618
rect 40910 39566 40962 39618
rect 51214 39566 51266 39618
rect 8318 39454 8370 39506
rect 17838 39454 17890 39506
rect 30382 39454 30434 39506
rect 41694 39454 41746 39506
rect 45614 39454 45666 39506
rect 53454 39454 53506 39506
rect 53678 39454 53730 39506
rect 10894 39342 10946 39394
rect 13806 39342 13858 39394
rect 20862 39342 20914 39394
rect 21534 39342 21586 39394
rect 37662 39342 37714 39394
rect 40014 39342 40066 39394
rect 46846 39342 46898 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 8542 39006 8594 39058
rect 10334 39006 10386 39058
rect 17950 39006 18002 39058
rect 26910 39006 26962 39058
rect 41918 39006 41970 39058
rect 43374 39006 43426 39058
rect 44046 39006 44098 39058
rect 47630 39006 47682 39058
rect 49646 39006 49698 39058
rect 51326 39006 51378 39058
rect 52334 39006 52386 39058
rect 5630 38894 5682 38946
rect 9886 38894 9938 38946
rect 11342 38894 11394 38946
rect 12238 38894 12290 38946
rect 13582 38894 13634 38946
rect 20974 38894 21026 38946
rect 25678 38894 25730 38946
rect 33630 38894 33682 38946
rect 40574 38894 40626 38946
rect 54014 38894 54066 38946
rect 4958 38782 5010 38834
rect 9774 38782 9826 38834
rect 10782 38782 10834 38834
rect 12798 38782 12850 38834
rect 20302 38782 20354 38834
rect 26798 38782 26850 38834
rect 27022 38782 27074 38834
rect 28366 38782 28418 38834
rect 31614 38782 31666 38834
rect 35086 38782 35138 38834
rect 42926 38782 42978 38834
rect 43150 38782 43202 38834
rect 43486 38782 43538 38834
rect 43934 38782 43986 38834
rect 44158 38782 44210 38834
rect 44606 38782 44658 38834
rect 47742 38782 47794 38834
rect 48414 38782 48466 38834
rect 49534 38782 49586 38834
rect 49758 38782 49810 38834
rect 51214 38782 51266 38834
rect 51662 38782 51714 38834
rect 53006 38782 53058 38834
rect 54350 38782 54402 38834
rect 7758 38670 7810 38722
rect 15710 38670 15762 38722
rect 23102 38670 23154 38722
rect 23550 38670 23602 38722
rect 29038 38670 29090 38722
rect 31166 38670 31218 38722
rect 36990 38670 37042 38722
rect 44382 38670 44434 38722
rect 48526 38670 48578 38722
rect 51438 38670 51490 38722
rect 53342 38670 53394 38722
rect 54126 38670 54178 38722
rect 27246 38558 27298 38610
rect 27470 38558 27522 38610
rect 47854 38558 47906 38610
rect 48750 38558 48802 38610
rect 49982 38558 50034 38610
rect 52894 38558 52946 38610
rect 53230 38558 53282 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 15710 38222 15762 38274
rect 52670 38222 52722 38274
rect 12686 38110 12738 38162
rect 25342 38110 25394 38162
rect 27470 38110 27522 38162
rect 32846 38110 32898 38162
rect 34974 38110 35026 38162
rect 36318 38110 36370 38162
rect 36654 38110 36706 38162
rect 37550 38110 37602 38162
rect 39678 38110 39730 38162
rect 41806 38110 41858 38162
rect 43934 38110 43986 38162
rect 47182 38110 47234 38162
rect 49310 38110 49362 38162
rect 52110 38110 52162 38162
rect 54238 38110 54290 38162
rect 56366 38110 56418 38162
rect 8318 37998 8370 38050
rect 15486 37998 15538 38050
rect 15934 37998 15986 38050
rect 16158 37998 16210 38050
rect 24558 37998 24610 38050
rect 32174 37998 32226 38050
rect 36430 37998 36482 38050
rect 40350 37998 40402 38050
rect 41022 37998 41074 38050
rect 49982 37998 50034 38050
rect 50654 37998 50706 38050
rect 52334 37998 52386 38050
rect 53454 37998 53506 38050
rect 8990 37886 9042 37938
rect 29598 37886 29650 37938
rect 30382 37886 30434 37938
rect 36766 37886 36818 37938
rect 50990 37886 51042 37938
rect 15598 37774 15650 37826
rect 27918 37774 27970 37826
rect 35534 37774 35586 37826
rect 44606 37774 44658 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 8766 37438 8818 37490
rect 11230 37438 11282 37490
rect 24222 37438 24274 37490
rect 38334 37438 38386 37490
rect 40686 37438 40738 37490
rect 41470 37438 41522 37490
rect 50094 37438 50146 37490
rect 10110 37326 10162 37378
rect 12574 37326 12626 37378
rect 15934 37326 15986 37378
rect 24894 37326 24946 37378
rect 27694 37326 27746 37378
rect 34638 37326 34690 37378
rect 37438 37326 37490 37378
rect 44942 37326 44994 37378
rect 52558 37326 52610 37378
rect 52670 37326 52722 37378
rect 52782 37326 52834 37378
rect 53454 37326 53506 37378
rect 53678 37326 53730 37378
rect 5406 37214 5458 37266
rect 11790 37214 11842 37266
rect 26686 37214 26738 37266
rect 31726 37214 31778 37266
rect 31950 37214 32002 37266
rect 33854 37214 33906 37266
rect 37326 37214 37378 37266
rect 37662 37214 37714 37266
rect 37886 37214 37938 37266
rect 45614 37214 45666 37266
rect 48190 37214 48242 37266
rect 48526 37214 48578 37266
rect 49534 37214 49586 37266
rect 49758 37214 49810 37266
rect 51102 37214 51154 37266
rect 51326 37214 51378 37266
rect 51550 37214 51602 37266
rect 53566 37214 53618 37266
rect 6190 37102 6242 37154
rect 8318 37102 8370 37154
rect 14702 37102 14754 37154
rect 17726 37102 17778 37154
rect 32510 37102 32562 37154
rect 36766 37102 36818 37154
rect 42366 37102 42418 37154
rect 42814 37102 42866 37154
rect 46174 37102 46226 37154
rect 52110 37102 52162 37154
rect 32174 36990 32226 37042
rect 32398 36990 32450 37042
rect 48078 36990 48130 37042
rect 48414 36990 48466 37042
rect 50990 36990 51042 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 7758 36654 7810 36706
rect 8654 36654 8706 36706
rect 7982 36542 8034 36594
rect 9102 36542 9154 36594
rect 11230 36542 11282 36594
rect 15262 36542 15314 36594
rect 17390 36542 17442 36594
rect 20862 36542 20914 36594
rect 25342 36542 25394 36594
rect 27470 36542 27522 36594
rect 27918 36542 27970 36594
rect 35310 36542 35362 36594
rect 37550 36542 37602 36594
rect 42254 36542 42306 36594
rect 48974 36542 49026 36594
rect 50542 36542 50594 36594
rect 52670 36542 52722 36594
rect 8206 36430 8258 36482
rect 12014 36430 12066 36482
rect 12462 36430 12514 36482
rect 14478 36430 14530 36482
rect 17950 36430 18002 36482
rect 24558 36430 24610 36482
rect 39454 36430 39506 36482
rect 42926 36430 42978 36482
rect 43150 36430 43202 36482
rect 43374 36430 43426 36482
rect 43598 36430 43650 36482
rect 46062 36430 46114 36482
rect 49870 36430 49922 36482
rect 6414 36318 6466 36370
rect 7534 36318 7586 36370
rect 18734 36318 18786 36370
rect 40126 36318 40178 36370
rect 46846 36318 46898 36370
rect 5742 36206 5794 36258
rect 13918 36206 13970 36258
rect 21982 36206 22034 36258
rect 29598 36206 29650 36258
rect 43038 36206 43090 36258
rect 44270 36206 44322 36258
rect 45502 36206 45554 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 19742 35870 19794 35922
rect 40350 35870 40402 35922
rect 41470 35870 41522 35922
rect 14030 35758 14082 35810
rect 18846 35758 18898 35810
rect 21870 35758 21922 35810
rect 29374 35758 29426 35810
rect 4510 35646 4562 35698
rect 7758 35646 7810 35698
rect 13246 35646 13298 35698
rect 16606 35646 16658 35698
rect 17614 35646 17666 35698
rect 21198 35646 21250 35698
rect 24446 35646 24498 35698
rect 28590 35646 28642 35698
rect 31950 35646 32002 35698
rect 43486 35646 43538 35698
rect 5182 35534 5234 35586
rect 7310 35534 7362 35586
rect 16158 35534 16210 35586
rect 23998 35534 24050 35586
rect 31502 35534 31554 35586
rect 36094 35534 36146 35586
rect 45390 35534 45442 35586
rect 48078 35534 48130 35586
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 22430 35086 22482 35138
rect 22990 35086 23042 35138
rect 23102 35086 23154 35138
rect 13694 34974 13746 35026
rect 16830 34974 16882 35026
rect 35870 34974 35922 35026
rect 40798 34974 40850 35026
rect 41806 34974 41858 35026
rect 43934 34974 43986 35026
rect 48974 34974 49026 35026
rect 14254 34862 14306 34914
rect 22542 34862 22594 34914
rect 22766 34862 22818 34914
rect 33070 34862 33122 34914
rect 37998 34862 38050 34914
rect 44718 34862 44770 34914
rect 46062 34862 46114 34914
rect 33742 34750 33794 34802
rect 38670 34750 38722 34802
rect 46846 34750 46898 34802
rect 24670 34638 24722 34690
rect 30158 34638 30210 34690
rect 36542 34638 36594 34690
rect 41358 34638 41410 34690
rect 45390 34638 45442 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 18286 34302 18338 34354
rect 32622 34302 32674 34354
rect 33854 34302 33906 34354
rect 38894 34302 38946 34354
rect 39454 34302 39506 34354
rect 47742 34302 47794 34354
rect 13694 34190 13746 34242
rect 17726 34190 17778 34242
rect 30046 34190 30098 34242
rect 37438 34190 37490 34242
rect 40798 34190 40850 34242
rect 6190 34078 6242 34130
rect 16718 34078 16770 34130
rect 18734 34078 18786 34130
rect 19630 34078 19682 34130
rect 29374 34078 29426 34130
rect 38222 34078 38274 34130
rect 41918 34078 41970 34130
rect 6862 33966 6914 34018
rect 8990 33966 9042 34018
rect 9774 33966 9826 34018
rect 20414 33966 20466 34018
rect 22542 33966 22594 34018
rect 22990 33966 23042 34018
rect 32174 33966 32226 34018
rect 35310 33966 35362 34018
rect 45390 33966 45442 34018
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 14366 33406 14418 33458
rect 16494 33406 16546 33458
rect 18622 33406 18674 33458
rect 20750 33406 20802 33458
rect 24446 33406 24498 33458
rect 26574 33406 26626 33458
rect 27806 33406 27858 33458
rect 32622 33406 32674 33458
rect 41246 33406 41298 33458
rect 43374 33406 43426 33458
rect 17166 33294 17218 33346
rect 17838 33294 17890 33346
rect 23774 33294 23826 33346
rect 36318 33294 36370 33346
rect 40574 33294 40626 33346
rect 7086 33182 7138 33234
rect 21646 33182 21698 33234
rect 11230 33070 11282 33122
rect 13694 33070 13746 33122
rect 22990 33070 23042 33122
rect 27246 33070 27298 33122
rect 36766 33070 36818 33122
rect 43822 33070 43874 33122
rect 45726 33070 45778 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 12238 32734 12290 32786
rect 16158 32734 16210 32786
rect 29598 32734 29650 32786
rect 13582 32622 13634 32674
rect 22766 32622 22818 32674
rect 28366 32622 28418 32674
rect 33630 32622 33682 32674
rect 36542 32622 36594 32674
rect 37998 32622 38050 32674
rect 46846 32622 46898 32674
rect 49870 32622 49922 32674
rect 12910 32510 12962 32562
rect 17838 32510 17890 32562
rect 21086 32510 21138 32562
rect 22094 32510 22146 32562
rect 29150 32510 29202 32562
rect 35870 32510 35922 32562
rect 36430 32510 36482 32562
rect 42814 32510 42866 32562
rect 15710 32398 15762 32450
rect 18510 32398 18562 32450
rect 20638 32398 20690 32450
rect 24894 32398 24946 32450
rect 26238 32398 26290 32450
rect 43598 32398 43650 32450
rect 45726 32398 45778 32450
rect 46174 32398 46226 32450
rect 35982 32286 36034 32338
rect 36206 32286 36258 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 10782 31838 10834 31890
rect 12910 31838 12962 31890
rect 16606 31838 16658 31890
rect 17166 31838 17218 31890
rect 19406 31838 19458 31890
rect 20862 31838 20914 31890
rect 26910 31838 26962 31890
rect 34750 31838 34802 31890
rect 38334 31838 38386 31890
rect 40462 31838 40514 31890
rect 10110 31726 10162 31778
rect 13806 31726 13858 31778
rect 24110 31726 24162 31778
rect 31950 31726 32002 31778
rect 32622 31726 32674 31778
rect 37550 31726 37602 31778
rect 46846 31726 46898 31778
rect 51214 31726 51266 31778
rect 14478 31614 14530 31666
rect 18286 31614 18338 31666
rect 24782 31614 24834 31666
rect 43822 31614 43874 31666
rect 49534 31614 49586 31666
rect 20302 31502 20354 31554
rect 21646 31502 21698 31554
rect 27358 31502 27410 31554
rect 35198 31502 35250 31554
rect 36766 31502 36818 31554
rect 40910 31502 40962 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 44942 31166 44994 31218
rect 6414 31054 6466 31106
rect 10110 31054 10162 31106
rect 21646 31054 21698 31106
rect 37886 31054 37938 31106
rect 46622 31054 46674 31106
rect 50318 31054 50370 31106
rect 5966 30942 6018 30994
rect 15038 30942 15090 30994
rect 15710 30942 15762 30994
rect 15934 30942 15986 30994
rect 16158 30942 16210 30994
rect 16270 30942 16322 30994
rect 18510 30942 18562 30994
rect 19070 30942 19122 30994
rect 26350 30942 26402 30994
rect 26798 30942 26850 30994
rect 27022 30942 27074 30994
rect 29710 30942 29762 30994
rect 33742 30942 33794 30994
rect 37102 30942 37154 30994
rect 41582 30942 41634 30994
rect 45950 30942 46002 30994
rect 49534 30942 49586 30994
rect 3054 30830 3106 30882
rect 5182 30830 5234 30882
rect 30382 30830 30434 30882
rect 32510 30830 32562 30882
rect 34414 30830 34466 30882
rect 36542 30830 36594 30882
rect 40014 30830 40066 30882
rect 40462 30830 40514 30882
rect 42366 30830 42418 30882
rect 44494 30830 44546 30882
rect 48750 30830 48802 30882
rect 52446 30830 52498 30882
rect 15598 30718 15650 30770
rect 26238 30718 26290 30770
rect 26574 30718 26626 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 20190 30382 20242 30434
rect 49310 30382 49362 30434
rect 49758 30382 49810 30434
rect 19182 30270 19234 30322
rect 20638 30270 20690 30322
rect 21646 30270 21698 30322
rect 32286 30270 32338 30322
rect 32734 30270 32786 30322
rect 33294 30270 33346 30322
rect 48526 30270 48578 30322
rect 49534 30270 49586 30322
rect 5854 30158 5906 30210
rect 6078 30158 6130 30210
rect 6302 30158 6354 30210
rect 15374 30158 15426 30210
rect 16382 30158 16434 30210
rect 20078 30158 20130 30210
rect 20414 30158 20466 30210
rect 38558 30158 38610 30210
rect 44158 30158 44210 30210
rect 45726 30158 45778 30210
rect 49086 30158 49138 30210
rect 13918 30046 13970 30098
rect 17054 30046 17106 30098
rect 20750 30046 20802 30098
rect 24782 30046 24834 30098
rect 30046 30046 30098 30098
rect 34078 30046 34130 30098
rect 40350 30046 40402 30098
rect 43486 30046 43538 30098
rect 46398 30046 46450 30098
rect 5966 29934 6018 29986
rect 23326 29934 23378 29986
rect 28142 29934 28194 29986
rect 30494 29934 30546 29986
rect 31726 29934 31778 29986
rect 49646 29934 49698 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 9662 29598 9714 29650
rect 13134 29598 13186 29650
rect 17726 29598 17778 29650
rect 40798 29598 40850 29650
rect 46510 29598 46562 29650
rect 5182 29486 5234 29538
rect 5406 29486 5458 29538
rect 11566 29486 11618 29538
rect 16942 29486 16994 29538
rect 19294 29486 19346 29538
rect 22766 29486 22818 29538
rect 27246 29486 27298 29538
rect 30718 29486 30770 29538
rect 8990 29374 9042 29426
rect 18622 29374 18674 29426
rect 21982 29374 22034 29426
rect 26574 29374 26626 29426
rect 29934 29374 29986 29426
rect 33742 29374 33794 29426
rect 36990 29374 37042 29426
rect 39454 29374 39506 29426
rect 39678 29374 39730 29426
rect 41582 29374 41634 29426
rect 45166 29374 45218 29426
rect 45614 29374 45666 29426
rect 49758 29374 49810 29426
rect 5518 29262 5570 29314
rect 6078 29262 6130 29314
rect 8206 29262 8258 29314
rect 21422 29262 21474 29314
rect 24894 29262 24946 29314
rect 29374 29262 29426 29314
rect 32846 29262 32898 29314
rect 34414 29262 34466 29314
rect 36542 29262 36594 29314
rect 39118 29262 39170 29314
rect 42366 29262 42418 29314
rect 44494 29262 44546 29314
rect 45390 29262 45442 29314
rect 45950 29262 46002 29314
rect 49534 29262 49586 29314
rect 39230 29150 39282 29202
rect 39790 29150 39842 29202
rect 45838 29150 45890 29202
rect 50094 29150 50146 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 6526 28814 6578 28866
rect 7534 28814 7586 28866
rect 25902 28814 25954 28866
rect 7422 28702 7474 28754
rect 10782 28702 10834 28754
rect 12910 28702 12962 28754
rect 17390 28702 17442 28754
rect 19518 28702 19570 28754
rect 20078 28702 20130 28754
rect 21758 28702 21810 28754
rect 34974 28702 35026 28754
rect 52670 28702 52722 28754
rect 5966 28590 6018 28642
rect 6190 28590 6242 28642
rect 9998 28590 10050 28642
rect 16718 28590 16770 28642
rect 25678 28590 25730 28642
rect 26126 28590 26178 28642
rect 26350 28590 26402 28642
rect 28254 28590 28306 28642
rect 30270 28590 30322 28642
rect 49758 28590 49810 28642
rect 7310 28478 7362 28530
rect 15710 28478 15762 28530
rect 42254 28478 42306 28530
rect 50542 28478 50594 28530
rect 13806 28366 13858 28418
rect 15150 28366 15202 28418
rect 15262 28366 15314 28418
rect 15486 28366 15538 28418
rect 25118 28366 25170 28418
rect 25790 28366 25842 28418
rect 28814 28366 28866 28418
rect 36318 28366 36370 28418
rect 38894 28366 38946 28418
rect 44270 28366 44322 28418
rect 49310 28366 49362 28418
rect 53342 28366 53394 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 21758 28030 21810 28082
rect 32062 28030 32114 28082
rect 34414 28030 34466 28082
rect 6078 27918 6130 27970
rect 6302 27918 6354 27970
rect 13694 27918 13746 27970
rect 20862 27918 20914 27970
rect 21198 27918 21250 27970
rect 22542 27918 22594 27970
rect 30494 27918 30546 27970
rect 36094 27918 36146 27970
rect 41582 27918 41634 27970
rect 44158 27918 44210 27970
rect 13022 27806 13074 27858
rect 20750 27806 20802 27858
rect 21534 27806 21586 27858
rect 25006 27806 25058 27858
rect 25678 27806 25730 27858
rect 31502 27806 31554 27858
rect 31726 27806 31778 27858
rect 32174 27806 32226 27858
rect 35310 27806 35362 27858
rect 43486 27806 43538 27858
rect 46734 27806 46786 27858
rect 48078 27806 48130 27858
rect 49534 27806 49586 27858
rect 15822 27694 15874 27746
rect 16382 27694 16434 27746
rect 38222 27694 38274 27746
rect 46286 27694 46338 27746
rect 48750 27694 48802 27746
rect 52110 27694 52162 27746
rect 6414 27582 6466 27634
rect 31950 27582 32002 27634
rect 48638 27582 48690 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 6526 27246 6578 27298
rect 14702 27246 14754 27298
rect 15038 27246 15090 27298
rect 6302 27134 6354 27186
rect 8990 27134 9042 27186
rect 9438 27134 9490 27186
rect 10782 27134 10834 27186
rect 12910 27134 12962 27186
rect 14814 27134 14866 27186
rect 25566 27134 25618 27186
rect 27694 27134 27746 27186
rect 32286 27134 32338 27186
rect 38670 27134 38722 27186
rect 40798 27134 40850 27186
rect 49310 27134 49362 27186
rect 52446 27134 52498 27186
rect 56702 27134 56754 27186
rect 8542 27022 8594 27074
rect 10110 27022 10162 27074
rect 15262 27022 15314 27074
rect 24894 27022 24946 27074
rect 35086 27022 35138 27074
rect 37886 27022 37938 27074
rect 41806 27022 41858 27074
rect 46510 27022 46562 27074
rect 49870 27022 49922 27074
rect 50094 27022 50146 27074
rect 50206 27022 50258 27074
rect 51662 27022 51714 27074
rect 53790 27022 53842 27074
rect 13582 26910 13634 26962
rect 20974 26910 21026 26962
rect 28142 26910 28194 26962
rect 34414 26910 34466 26962
rect 41694 26910 41746 26962
rect 41918 26910 41970 26962
rect 47182 26910 47234 26962
rect 51214 26910 51266 26962
rect 51550 26910 51602 26962
rect 52334 26910 52386 26962
rect 54574 26910 54626 26962
rect 6862 26798 6914 26850
rect 8206 26798 8258 26850
rect 15150 26798 15202 26850
rect 18286 26798 18338 26850
rect 23214 26798 23266 26850
rect 42366 26798 42418 26850
rect 50654 26798 50706 26850
rect 51326 26798 51378 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 8878 26462 8930 26514
rect 11454 26462 11506 26514
rect 24894 26462 24946 26514
rect 31838 26462 31890 26514
rect 33742 26462 33794 26514
rect 42142 26462 42194 26514
rect 48414 26462 48466 26514
rect 49758 26462 49810 26514
rect 53230 26462 53282 26514
rect 54014 26462 54066 26514
rect 9998 26350 10050 26402
rect 18510 26350 18562 26402
rect 22318 26350 22370 26402
rect 29262 26350 29314 26402
rect 32398 26350 32450 26402
rect 35758 26350 35810 26402
rect 49870 26350 49922 26402
rect 49982 26350 50034 26402
rect 51326 26350 51378 26402
rect 53678 26350 53730 26402
rect 3390 26238 3442 26290
rect 7310 26238 7362 26290
rect 7534 26238 7586 26290
rect 8542 26238 8594 26290
rect 8990 26238 9042 26290
rect 9886 26238 9938 26290
rect 17838 26238 17890 26290
rect 21646 26238 21698 26290
rect 28590 26238 28642 26290
rect 40238 26238 40290 26290
rect 41582 26238 41634 26290
rect 42254 26238 42306 26290
rect 43598 26238 43650 26290
rect 48078 26238 48130 26290
rect 48414 26238 48466 26290
rect 48750 26238 48802 26290
rect 49534 26238 49586 26290
rect 51438 26238 51490 26290
rect 56142 26238 56194 26290
rect 4174 26126 4226 26178
rect 6302 26126 6354 26178
rect 6862 26126 6914 26178
rect 20638 26126 20690 26178
rect 24446 26126 24498 26178
rect 31390 26126 31442 26178
rect 42030 26126 42082 26178
rect 42814 26126 42866 26178
rect 44270 26126 44322 26178
rect 46398 26126 46450 26178
rect 46846 26126 46898 26178
rect 47518 26126 47570 26178
rect 49870 26126 49922 26178
rect 55358 26126 55410 26178
rect 7870 26014 7922 26066
rect 8766 26014 8818 26066
rect 9774 26014 9826 26066
rect 41806 26014 41858 26066
rect 42590 26014 42642 26066
rect 42926 26014 42978 26066
rect 51326 26014 51378 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 6190 25678 6242 25730
rect 6302 25678 6354 25730
rect 6526 25678 6578 25730
rect 6638 25678 6690 25730
rect 20526 25678 20578 25730
rect 20862 25678 20914 25730
rect 44382 25678 44434 25730
rect 50094 25678 50146 25730
rect 7870 25566 7922 25618
rect 9998 25566 10050 25618
rect 11230 25566 11282 25618
rect 18622 25566 18674 25618
rect 20302 25566 20354 25618
rect 22990 25566 23042 25618
rect 25118 25566 25170 25618
rect 25566 25566 25618 25618
rect 32174 25566 32226 25618
rect 34302 25566 34354 25618
rect 40798 25566 40850 25618
rect 42926 25566 42978 25618
rect 45838 25566 45890 25618
rect 50430 25566 50482 25618
rect 10782 25454 10834 25506
rect 15822 25454 15874 25506
rect 20190 25454 20242 25506
rect 20750 25454 20802 25506
rect 22318 25454 22370 25506
rect 31390 25454 31442 25506
rect 34750 25454 34802 25506
rect 40126 25454 40178 25506
rect 45950 25454 46002 25506
rect 48750 25454 48802 25506
rect 49758 25454 49810 25506
rect 51102 25454 51154 25506
rect 51550 25454 51602 25506
rect 52446 25454 52498 25506
rect 16494 25342 16546 25394
rect 37662 25342 37714 25394
rect 44718 25342 44770 25394
rect 45502 25342 45554 25394
rect 49534 25342 49586 25394
rect 49982 25342 50034 25394
rect 50878 25342 50930 25394
rect 51214 25342 51266 25394
rect 13694 25230 13746 25282
rect 19518 25230 19570 25282
rect 28254 25230 28306 25282
rect 38222 25230 38274 25282
rect 43374 25230 43426 25282
rect 44494 25230 44546 25282
rect 48414 25230 48466 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 17726 24894 17778 24946
rect 44942 24894 44994 24946
rect 48862 24894 48914 24946
rect 6974 24782 7026 24834
rect 14926 24782 14978 24834
rect 19630 24782 19682 24834
rect 25678 24782 25730 24834
rect 28142 24782 28194 24834
rect 36990 24782 37042 24834
rect 39678 24782 39730 24834
rect 45502 24782 45554 24834
rect 49534 24782 49586 24834
rect 49870 24782 49922 24834
rect 7310 24670 7362 24722
rect 13022 24670 13074 24722
rect 18846 24670 18898 24722
rect 27470 24670 27522 24722
rect 36206 24670 36258 24722
rect 45838 24670 45890 24722
rect 51214 24670 51266 24722
rect 55358 24670 55410 24722
rect 7086 24558 7138 24610
rect 18286 24558 18338 24610
rect 21758 24558 21810 24610
rect 22206 24558 22258 24610
rect 30270 24558 30322 24610
rect 39118 24558 39170 24610
rect 45614 24558 45666 24610
rect 51438 24558 51490 24610
rect 51886 24558 51938 24610
rect 52446 24558 52498 24610
rect 54574 24558 54626 24610
rect 55918 24558 55970 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 30046 24110 30098 24162
rect 34414 24110 34466 24162
rect 34638 24110 34690 24162
rect 52334 24110 52386 24162
rect 52670 24110 52722 24162
rect 12238 23998 12290 24050
rect 16606 23998 16658 24050
rect 17054 23998 17106 24050
rect 24670 23998 24722 24050
rect 26798 23998 26850 24050
rect 28030 23998 28082 24050
rect 29710 23998 29762 24050
rect 38334 23998 38386 24050
rect 40462 23998 40514 24050
rect 42590 23998 42642 24050
rect 44718 23998 44770 24050
rect 51326 23998 51378 24050
rect 9438 23886 9490 23938
rect 13694 23886 13746 23938
rect 23998 23886 24050 23938
rect 29822 23886 29874 23938
rect 30270 23886 30322 23938
rect 31390 23886 31442 23938
rect 31726 23886 31778 23938
rect 32174 23886 32226 23938
rect 34302 23886 34354 23938
rect 34862 23886 34914 23938
rect 34974 23886 35026 23938
rect 37550 23886 37602 23938
rect 41806 23886 41858 23938
rect 47070 23886 47122 23938
rect 48302 23886 48354 23938
rect 51662 23886 51714 23938
rect 10110 23774 10162 23826
rect 12910 23774 12962 23826
rect 14478 23774 14530 23826
rect 30382 23774 30434 23826
rect 31502 23774 31554 23826
rect 45614 23774 45666 23826
rect 45726 23774 45778 23826
rect 45838 23774 45890 23826
rect 51102 23774 51154 23826
rect 4622 23662 4674 23714
rect 5742 23662 5794 23714
rect 18958 23662 19010 23714
rect 27358 23662 27410 23714
rect 28478 23662 28530 23714
rect 32398 23662 32450 23714
rect 32846 23662 32898 23714
rect 41022 23662 41074 23714
rect 46286 23662 46338 23714
rect 46846 23662 46898 23714
rect 48078 23662 48130 23714
rect 51326 23662 51378 23714
rect 52558 23662 52610 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 10334 23326 10386 23378
rect 11230 23326 11282 23378
rect 16606 23326 16658 23378
rect 26350 23326 26402 23378
rect 48526 23326 48578 23378
rect 51214 23326 51266 23378
rect 3390 23214 3442 23266
rect 9662 23214 9714 23266
rect 13358 23214 13410 23266
rect 16046 23214 16098 23266
rect 20190 23214 20242 23266
rect 23438 23214 23490 23266
rect 38670 23214 38722 23266
rect 44942 23214 44994 23266
rect 2718 23102 2770 23154
rect 6078 23102 6130 23154
rect 12014 23102 12066 23154
rect 12686 23102 12738 23154
rect 19182 23102 19234 23154
rect 26910 23102 26962 23154
rect 36542 23102 36594 23154
rect 37998 23102 38050 23154
rect 42030 23102 42082 23154
rect 48750 23102 48802 23154
rect 49534 23102 49586 23154
rect 49758 23102 49810 23154
rect 50430 23102 50482 23154
rect 52222 23102 52274 23154
rect 52558 23102 52610 23154
rect 52782 23102 52834 23154
rect 5518 22990 5570 23042
rect 6862 22990 6914 23042
rect 8990 22990 9042 23042
rect 15486 22990 15538 23042
rect 28926 22990 28978 23042
rect 33630 22990 33682 23042
rect 35758 22990 35810 23042
rect 40798 22990 40850 23042
rect 47294 22990 47346 23042
rect 48638 22990 48690 23042
rect 51774 22990 51826 23042
rect 52446 22990 52498 23042
rect 51550 22878 51602 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 12350 22542 12402 22594
rect 12574 22542 12626 22594
rect 41582 22542 41634 22594
rect 41918 22542 41970 22594
rect 47182 22542 47234 22594
rect 47742 22542 47794 22594
rect 51662 22542 51714 22594
rect 1822 22430 1874 22482
rect 3950 22430 4002 22482
rect 8430 22430 8482 22482
rect 13582 22430 13634 22482
rect 15262 22430 15314 22482
rect 17390 22430 17442 22482
rect 18734 22430 18786 22482
rect 20862 22430 20914 22482
rect 24558 22430 24610 22482
rect 26686 22430 26738 22482
rect 28814 22430 28866 22482
rect 31838 22430 31890 22482
rect 33966 22430 34018 22482
rect 35086 22430 35138 22482
rect 38670 22430 38722 22482
rect 40798 22430 40850 22482
rect 4734 22318 4786 22370
rect 6638 22318 6690 22370
rect 12014 22318 12066 22370
rect 12126 22318 12178 22370
rect 14590 22318 14642 22370
rect 17950 22318 18002 22370
rect 21646 22318 21698 22370
rect 26014 22318 26066 22370
rect 31166 22318 31218 22370
rect 37998 22318 38050 22370
rect 41358 22318 41410 22370
rect 41806 22318 41858 22370
rect 46174 22318 46226 22370
rect 46958 22318 47010 22370
rect 47966 22318 48018 22370
rect 48078 22318 48130 22370
rect 51214 22318 51266 22370
rect 51438 22318 51490 22370
rect 51998 22318 52050 22370
rect 12686 22206 12738 22258
rect 22430 22206 22482 22258
rect 34638 22206 34690 22258
rect 46286 22206 46338 22258
rect 46510 22206 46562 22258
rect 47630 22206 47682 22258
rect 42366 22094 42418 22146
rect 51998 22094 52050 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 4958 21758 5010 21810
rect 7310 21758 7362 21810
rect 13134 21758 13186 21810
rect 14142 21758 14194 21810
rect 20862 21758 20914 21810
rect 21310 21758 21362 21810
rect 22318 21758 22370 21810
rect 23998 21758 24050 21810
rect 46062 21758 46114 21810
rect 50878 21758 50930 21810
rect 25678 21646 25730 21698
rect 28366 21646 28418 21698
rect 35646 21646 35698 21698
rect 41470 21646 41522 21698
rect 45614 21646 45666 21698
rect 45838 21646 45890 21698
rect 46398 21646 46450 21698
rect 46846 21646 46898 21698
rect 55358 21646 55410 21698
rect 1822 21534 1874 21586
rect 9886 21534 9938 21586
rect 24110 21534 24162 21586
rect 27694 21534 27746 21586
rect 34974 21534 35026 21586
rect 39342 21534 39394 21586
rect 42142 21534 42194 21586
rect 46286 21534 46338 21586
rect 46846 21534 46898 21586
rect 47070 21534 47122 21586
rect 47294 21534 47346 21586
rect 51438 21534 51490 21586
rect 2494 21422 2546 21474
rect 10558 21422 10610 21474
rect 12686 21422 12738 21474
rect 30494 21422 30546 21474
rect 42926 21422 42978 21474
rect 45054 21422 45106 21474
rect 23998 21310 24050 21362
rect 24334 21310 24386 21362
rect 24558 21310 24610 21362
rect 47406 21310 47458 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 5630 20862 5682 20914
rect 11902 20862 11954 20914
rect 20862 20862 20914 20914
rect 23214 20862 23266 20914
rect 25342 20862 25394 20914
rect 28814 20862 28866 20914
rect 32510 20862 32562 20914
rect 32958 20862 33010 20914
rect 36542 20862 36594 20914
rect 42142 20862 42194 20914
rect 45390 20862 45442 20914
rect 46174 20862 46226 20914
rect 48750 20862 48802 20914
rect 50878 20862 50930 20914
rect 9102 20750 9154 20802
rect 17950 20750 18002 20802
rect 22542 20750 22594 20802
rect 26014 20750 26066 20802
rect 29710 20750 29762 20802
rect 33742 20750 33794 20802
rect 39230 20750 39282 20802
rect 45950 20750 46002 20802
rect 48078 20750 48130 20802
rect 9774 20638 9826 20690
rect 18734 20638 18786 20690
rect 26686 20638 26738 20690
rect 30382 20638 30434 20690
rect 34414 20638 34466 20690
rect 40014 20638 40066 20690
rect 46286 20638 46338 20690
rect 3166 20526 3218 20578
rect 3838 20526 3890 20578
rect 6526 20526 6578 20578
rect 12350 20526 12402 20578
rect 14814 20526 14866 20578
rect 15486 20526 15538 20578
rect 17054 20526 17106 20578
rect 21870 20526 21922 20578
rect 37550 20526 37602 20578
rect 38110 20526 38162 20578
rect 38558 20526 38610 20578
rect 42590 20526 42642 20578
rect 51326 20526 51378 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 9886 20190 9938 20242
rect 10670 20190 10722 20242
rect 19518 20190 19570 20242
rect 20638 20190 20690 20242
rect 27470 20190 27522 20242
rect 29822 20190 29874 20242
rect 34302 20190 34354 20242
rect 38558 20190 38610 20242
rect 40574 20190 40626 20242
rect 50542 20190 50594 20242
rect 54910 20190 54962 20242
rect 2942 20078 2994 20130
rect 6414 20078 6466 20130
rect 8990 20078 9042 20130
rect 14702 20078 14754 20130
rect 21982 20078 22034 20130
rect 31166 20078 31218 20130
rect 35646 20078 35698 20130
rect 38446 20078 38498 20130
rect 39902 20078 39954 20130
rect 43710 20078 43762 20130
rect 47294 20078 47346 20130
rect 49982 20078 50034 20130
rect 53678 20078 53730 20130
rect 2158 19966 2210 20018
rect 5630 19966 5682 20018
rect 14030 19966 14082 20018
rect 18062 19966 18114 20018
rect 18510 19966 18562 20018
rect 21198 19966 21250 20018
rect 30942 19966 30994 20018
rect 34862 19966 34914 20018
rect 38334 19966 38386 20018
rect 39342 19966 39394 20018
rect 48078 19966 48130 20018
rect 54462 19966 54514 20018
rect 5070 19854 5122 19906
rect 8542 19854 8594 19906
rect 16830 19854 16882 19906
rect 18286 19854 18338 19906
rect 24110 19854 24162 19906
rect 24558 19854 24610 19906
rect 25566 19854 25618 19906
rect 31278 19854 31330 19906
rect 37774 19854 37826 19906
rect 45166 19854 45218 19906
rect 48526 19854 48578 19906
rect 51550 19854 51602 19906
rect 17726 19742 17778 19794
rect 17838 19742 17890 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 6302 19406 6354 19458
rect 6526 19406 6578 19458
rect 6750 19406 6802 19458
rect 2830 19294 2882 19346
rect 4958 19294 5010 19346
rect 6078 19294 6130 19346
rect 12574 19294 12626 19346
rect 13582 19294 13634 19346
rect 21534 19294 21586 19346
rect 22990 19294 23042 19346
rect 33518 19294 33570 19346
rect 40910 19294 40962 19346
rect 41358 19294 41410 19346
rect 49646 19294 49698 19346
rect 51774 19294 51826 19346
rect 53454 19294 53506 19346
rect 2158 19182 2210 19234
rect 9662 19182 9714 19234
rect 15598 19182 15650 19234
rect 23550 19182 23602 19234
rect 30606 19182 30658 19234
rect 38110 19182 38162 19234
rect 48862 19182 48914 19234
rect 56254 19182 56306 19234
rect 56814 19182 56866 19234
rect 10446 19070 10498 19122
rect 20078 19070 20130 19122
rect 25566 19070 25618 19122
rect 31390 19070 31442 19122
rect 38782 19070 38834 19122
rect 52670 19070 52722 19122
rect 55582 19070 55634 19122
rect 7198 18958 7250 19010
rect 33966 18958 34018 19010
rect 46510 18958 46562 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 5294 18622 5346 18674
rect 10670 18622 10722 18674
rect 31614 18622 31666 18674
rect 38894 18622 38946 18674
rect 53678 18622 53730 18674
rect 13246 18510 13298 18562
rect 23662 18510 23714 18562
rect 43934 18510 43986 18562
rect 54798 18510 54850 18562
rect 7646 18398 7698 18450
rect 7870 18398 7922 18450
rect 8206 18398 8258 18450
rect 13134 18398 13186 18450
rect 13470 18398 13522 18450
rect 14142 18398 14194 18450
rect 17950 18398 18002 18450
rect 21310 18398 21362 18450
rect 21758 18398 21810 18450
rect 25678 18398 25730 18450
rect 34078 18398 34130 18450
rect 37438 18398 37490 18450
rect 40798 18398 40850 18450
rect 41918 18398 41970 18450
rect 49646 18398 49698 18450
rect 50318 18398 50370 18450
rect 53342 18398 53394 18450
rect 53566 18398 53618 18450
rect 14814 18286 14866 18338
rect 16942 18286 16994 18338
rect 18622 18286 18674 18338
rect 20750 18286 20802 18338
rect 21982 18286 22034 18338
rect 26462 18286 26514 18338
rect 28590 18286 28642 18338
rect 29038 18286 29090 18338
rect 34862 18286 34914 18338
rect 36990 18286 37042 18338
rect 52446 18286 52498 18338
rect 8430 18174 8482 18226
rect 12686 18174 12738 18226
rect 22206 18174 22258 18226
rect 22430 18174 22482 18226
rect 22542 18174 22594 18226
rect 53230 18174 53282 18226
rect 53790 18174 53842 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 12686 17726 12738 17778
rect 13582 17726 13634 17778
rect 17278 17726 17330 17778
rect 22654 17726 22706 17778
rect 24782 17726 24834 17778
rect 44494 17726 44546 17778
rect 45502 17726 45554 17778
rect 47630 17726 47682 17778
rect 53790 17726 53842 17778
rect 55918 17726 55970 17778
rect 57150 17726 57202 17778
rect 8318 17614 8370 17666
rect 25454 17614 25506 17666
rect 41694 17614 41746 17666
rect 48302 17614 48354 17666
rect 56702 17614 56754 17666
rect 18846 17502 18898 17554
rect 26462 17502 26514 17554
rect 35086 17502 35138 17554
rect 41022 17502 41074 17554
rect 42366 17502 42418 17554
rect 6526 17390 6578 17442
rect 20190 17390 20242 17442
rect 29598 17390 29650 17442
rect 48862 17390 48914 17442
rect 51998 17390 52050 17442
rect 52670 17390 52722 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 22654 17054 22706 17106
rect 25790 17054 25842 17106
rect 27582 17054 27634 17106
rect 34750 17054 34802 17106
rect 36766 17054 36818 17106
rect 48750 17054 48802 17106
rect 6414 16942 6466 16994
rect 9774 16942 9826 16994
rect 14926 16942 14978 16994
rect 17726 16942 17778 16994
rect 20078 16942 20130 16994
rect 31614 16942 31666 16994
rect 33742 16942 33794 16994
rect 35198 16942 35250 16994
rect 37326 16942 37378 16994
rect 39790 16942 39842 16994
rect 43486 16942 43538 16994
rect 51550 16942 51602 16994
rect 5070 16830 5122 16882
rect 5742 16830 5794 16882
rect 8990 16830 9042 16882
rect 10782 16830 10834 16882
rect 11454 16830 11506 16882
rect 19406 16830 19458 16882
rect 23326 16830 23378 16882
rect 28142 16830 28194 16882
rect 28926 16830 28978 16882
rect 33630 16830 33682 16882
rect 34638 16830 34690 16882
rect 37550 16830 37602 16882
rect 38222 16830 38274 16882
rect 38558 16830 38610 16882
rect 42814 16830 42866 16882
rect 46062 16830 46114 16882
rect 49534 16830 49586 16882
rect 2158 16718 2210 16770
rect 4286 16718 4338 16770
rect 8542 16718 8594 16770
rect 12126 16718 12178 16770
rect 14254 16718 14306 16770
rect 22206 16718 22258 16770
rect 23550 16718 23602 16770
rect 31054 16718 31106 16770
rect 45614 16718 45666 16770
rect 48302 16718 48354 16770
rect 23886 16606 23938 16658
rect 38558 16606 38610 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 13918 16270 13970 16322
rect 14142 16270 14194 16322
rect 37662 16270 37714 16322
rect 37998 16270 38050 16322
rect 5630 16158 5682 16210
rect 9438 16158 9490 16210
rect 11566 16158 11618 16210
rect 12798 16158 12850 16210
rect 13806 16158 13858 16210
rect 17278 16158 17330 16210
rect 19406 16158 19458 16210
rect 19854 16158 19906 16210
rect 30830 16158 30882 16210
rect 32958 16158 33010 16210
rect 37774 16158 37826 16210
rect 38782 16158 38834 16210
rect 40910 16158 40962 16210
rect 45502 16158 45554 16210
rect 52670 16158 52722 16210
rect 8766 16046 8818 16098
rect 14366 16046 14418 16098
rect 16606 16046 16658 16098
rect 30046 16046 30098 16098
rect 38222 16046 38274 16098
rect 41694 16046 41746 16098
rect 48302 16046 48354 16098
rect 49758 16046 49810 16098
rect 4510 15934 4562 15986
rect 12238 15934 12290 15986
rect 44046 15934 44098 15986
rect 47630 15934 47682 15986
rect 50542 15934 50594 15986
rect 53454 15934 53506 15986
rect 13806 15822 13858 15874
rect 23774 15822 23826 15874
rect 27134 15822 27186 15874
rect 33518 15822 33570 15874
rect 34078 15822 34130 15874
rect 36430 15822 36482 15874
rect 42142 15822 42194 15874
rect 44718 15822 44770 15874
rect 49198 15822 49250 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 38894 15486 38946 15538
rect 52894 15486 52946 15538
rect 53342 15486 53394 15538
rect 15262 15374 15314 15426
rect 26910 15374 26962 15426
rect 36318 15374 36370 15426
rect 42254 15374 42306 15426
rect 48414 15374 48466 15426
rect 50318 15374 50370 15426
rect 54126 15374 54178 15426
rect 16046 15262 16098 15314
rect 18846 15262 18898 15314
rect 19518 15262 19570 15314
rect 26238 15262 26290 15314
rect 35646 15262 35698 15314
rect 45614 15262 45666 15314
rect 45838 15262 45890 15314
rect 46062 15262 46114 15314
rect 46286 15262 46338 15314
rect 49646 15262 49698 15314
rect 10110 15150 10162 15202
rect 13134 15150 13186 15202
rect 16606 15150 16658 15202
rect 21534 15150 21586 15202
rect 29038 15150 29090 15202
rect 38446 15150 38498 15202
rect 52446 15150 52498 15202
rect 9998 15038 10050 15090
rect 46398 15038 46450 15090
rect 52670 15038 52722 15090
rect 53342 15038 53394 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 10782 14590 10834 14642
rect 11342 14590 11394 14642
rect 19742 14590 19794 14642
rect 20190 14590 20242 14642
rect 22542 14590 22594 14642
rect 24670 14590 24722 14642
rect 28142 14590 28194 14642
rect 32734 14590 32786 14642
rect 34862 14590 34914 14642
rect 41694 14590 41746 14642
rect 43822 14590 43874 14642
rect 48190 14590 48242 14642
rect 50318 14590 50370 14642
rect 50766 14590 50818 14642
rect 53454 14590 53506 14642
rect 55582 14590 55634 14642
rect 7982 14478 8034 14530
rect 16830 14478 16882 14530
rect 21758 14478 21810 14530
rect 25342 14478 25394 14530
rect 32062 14478 32114 14530
rect 39566 14478 39618 14530
rect 47518 14478 47570 14530
rect 56366 14478 56418 14530
rect 56814 14478 56866 14530
rect 8654 14366 8706 14418
rect 17614 14366 17666 14418
rect 26014 14366 26066 14418
rect 16270 14254 16322 14306
rect 20862 14254 20914 14306
rect 30046 14254 30098 14306
rect 30942 14254 30994 14306
rect 35310 14254 35362 14306
rect 36318 14254 36370 14306
rect 46286 14254 46338 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 17838 13918 17890 13970
rect 23886 13918 23938 13970
rect 26014 13918 26066 13970
rect 33518 13918 33570 13970
rect 38782 13918 38834 13970
rect 53678 13918 53730 13970
rect 6974 13806 7026 13858
rect 8094 13806 8146 13858
rect 8654 13806 8706 13858
rect 21310 13806 21362 13858
rect 36206 13806 36258 13858
rect 40014 13806 40066 13858
rect 3502 13694 3554 13746
rect 8990 13694 9042 13746
rect 9998 13694 10050 13746
rect 10446 13694 10498 13746
rect 10894 13694 10946 13746
rect 14030 13694 14082 13746
rect 20638 13694 20690 13746
rect 26910 13694 26962 13746
rect 35534 13694 35586 13746
rect 46958 13694 47010 13746
rect 47854 13694 47906 13746
rect 53118 13694 53170 13746
rect 53342 13694 53394 13746
rect 53566 13694 53618 13746
rect 53790 13694 53842 13746
rect 4174 13582 4226 13634
rect 6302 13582 6354 13634
rect 6862 13582 6914 13634
rect 7758 13582 7810 13634
rect 10222 13582 10274 13634
rect 11118 13582 11170 13634
rect 14814 13582 14866 13634
rect 16942 13582 16994 13634
rect 23438 13582 23490 13634
rect 29150 13582 29202 13634
rect 38334 13582 38386 13634
rect 45390 13582 45442 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19294 13134 19346 13186
rect 19518 13134 19570 13186
rect 27918 13134 27970 13186
rect 28030 13134 28082 13186
rect 28254 13134 28306 13186
rect 28478 13134 28530 13186
rect 6974 13022 7026 13074
rect 19070 13022 19122 13074
rect 19966 13022 20018 13074
rect 23326 13022 23378 13074
rect 30718 13022 30770 13074
rect 32846 13022 32898 13074
rect 33406 13022 33458 13074
rect 39790 13022 39842 13074
rect 41918 13022 41970 13074
rect 48414 13022 48466 13074
rect 6078 12910 6130 12962
rect 7086 12910 7138 12962
rect 8990 12910 9042 12962
rect 9550 12910 9602 12962
rect 10670 12910 10722 12962
rect 11006 12910 11058 12962
rect 12574 12910 12626 12962
rect 12798 12910 12850 12962
rect 23214 12910 23266 12962
rect 23550 12910 23602 12962
rect 29934 12910 29986 12962
rect 36318 12910 36370 12962
rect 39118 12910 39170 12962
rect 45502 12910 45554 12962
rect 53454 12910 53506 12962
rect 53678 12910 53730 12962
rect 6638 12798 6690 12850
rect 9102 12798 9154 12850
rect 11342 12798 11394 12850
rect 11902 12798 11954 12850
rect 15598 12798 15650 12850
rect 18846 12798 18898 12850
rect 28590 12798 28642 12850
rect 35534 12798 35586 12850
rect 44046 12798 44098 12850
rect 46286 12798 46338 12850
rect 54126 12798 54178 12850
rect 5742 12686 5794 12738
rect 6862 12686 6914 12738
rect 7198 12686 7250 12738
rect 7758 12686 7810 12738
rect 9214 12686 9266 12738
rect 11006 12686 11058 12738
rect 14030 12686 14082 12738
rect 16718 12686 16770 12738
rect 17278 12686 17330 12738
rect 21646 12686 21698 12738
rect 23886 12686 23938 12738
rect 26350 12686 26402 12738
rect 36766 12686 36818 12738
rect 48862 12686 48914 12738
rect 53342 12686 53394 12738
rect 53902 12686 53954 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 9774 12350 9826 12402
rect 23886 12350 23938 12402
rect 33966 12350 34018 12402
rect 40238 12350 40290 12402
rect 54462 12350 54514 12402
rect 55022 12350 55074 12402
rect 10334 12238 10386 12290
rect 11678 12238 11730 12290
rect 14366 12238 14418 12290
rect 20750 12238 20802 12290
rect 24334 12238 24386 12290
rect 29934 12238 29986 12290
rect 42366 12238 42418 12290
rect 47630 12238 47682 12290
rect 49534 12238 49586 12290
rect 8990 12126 9042 12178
rect 11006 12126 11058 12178
rect 14478 12126 14530 12178
rect 15262 12126 15314 12178
rect 15598 12126 15650 12178
rect 19966 12126 20018 12178
rect 24110 12126 24162 12178
rect 26686 12126 26738 12178
rect 28030 12126 28082 12178
rect 28590 12126 28642 12178
rect 29150 12126 29202 12178
rect 36990 12126 37042 12178
rect 41582 12126 41634 12178
rect 48414 12126 48466 12178
rect 53678 12126 53730 12178
rect 3950 12014 4002 12066
rect 13806 12014 13858 12066
rect 22878 12014 22930 12066
rect 23438 12014 23490 12066
rect 26126 12014 26178 12066
rect 32062 12014 32114 12066
rect 37662 12014 37714 12066
rect 39790 12014 39842 12066
rect 44494 12014 44546 12066
rect 45502 12014 45554 12066
rect 50766 12014 50818 12066
rect 52894 12014 52946 12066
rect 10110 11902 10162 11954
rect 14254 11902 14306 11954
rect 24222 11902 24274 11954
rect 26126 11902 26178 11954
rect 26462 11902 26514 11954
rect 26686 11902 26738 11954
rect 27022 11902 27074 11954
rect 28366 11902 28418 11954
rect 54238 11902 54290 11954
rect 54574 11902 54626 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 12798 11566 12850 11618
rect 25006 11566 25058 11618
rect 38334 11566 38386 11618
rect 45726 11566 45778 11618
rect 45838 11566 45890 11618
rect 46062 11566 46114 11618
rect 52334 11566 52386 11618
rect 53566 11566 53618 11618
rect 54238 11566 54290 11618
rect 8654 11454 8706 11506
rect 20414 11454 20466 11506
rect 28366 11454 28418 11506
rect 31950 11454 32002 11506
rect 36206 11454 36258 11506
rect 38446 11454 38498 11506
rect 39118 11454 39170 11506
rect 48862 11454 48914 11506
rect 50990 11454 51042 11506
rect 53678 11454 53730 11506
rect 5742 11342 5794 11394
rect 9998 11342 10050 11394
rect 13022 11342 13074 11394
rect 16158 11342 16210 11394
rect 21982 11342 22034 11394
rect 23550 11342 23602 11394
rect 24222 11342 24274 11394
rect 24670 11342 24722 11394
rect 25566 11342 25618 11394
rect 35758 11342 35810 11394
rect 46286 11342 46338 11394
rect 46846 11342 46898 11394
rect 47518 11342 47570 11394
rect 48190 11342 48242 11394
rect 51998 11342 52050 11394
rect 53902 11342 53954 11394
rect 54126 11342 54178 11394
rect 6526 11230 6578 11282
rect 10222 11230 10274 11282
rect 16830 11230 16882 11282
rect 22318 11230 22370 11282
rect 23662 11230 23714 11282
rect 26238 11230 26290 11282
rect 46398 11230 46450 11282
rect 47406 11230 47458 11282
rect 52222 11230 52274 11282
rect 9214 11118 9266 11170
rect 10670 11118 10722 11170
rect 11902 11118 11954 11170
rect 12462 11118 12514 11170
rect 12686 11118 12738 11170
rect 14030 11118 14082 11170
rect 22206 11118 22258 11170
rect 38558 11118 38610 11170
rect 47182 11118 47234 11170
rect 51438 11118 51490 11170
rect 54910 11118 54962 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 6750 10782 6802 10834
rect 10110 10782 10162 10834
rect 12238 10782 12290 10834
rect 12798 10782 12850 10834
rect 32174 10782 32226 10834
rect 40014 10782 40066 10834
rect 10670 10670 10722 10722
rect 12126 10670 12178 10722
rect 16718 10670 16770 10722
rect 22878 10670 22930 10722
rect 27022 10670 27074 10722
rect 39454 10670 39506 10722
rect 41806 10670 41858 10722
rect 42814 10670 42866 10722
rect 45950 10670 46002 10722
rect 46622 10670 46674 10722
rect 48638 10670 48690 10722
rect 56366 10670 56418 10722
rect 2830 10558 2882 10610
rect 3166 10558 3218 10610
rect 3390 10558 3442 10610
rect 4398 10558 4450 10610
rect 6638 10558 6690 10610
rect 6974 10558 7026 10610
rect 7422 10558 7474 10610
rect 9774 10558 9826 10610
rect 11006 10558 11058 10610
rect 19070 10558 19122 10610
rect 22430 10558 22482 10610
rect 22654 10558 22706 10610
rect 27918 10558 27970 10610
rect 32286 10558 32338 10610
rect 32510 10558 32562 10610
rect 32734 10558 32786 10610
rect 38446 10558 38498 10610
rect 39342 10558 39394 10610
rect 45166 10558 45218 10610
rect 51438 10558 51490 10610
rect 3054 10446 3106 10498
rect 3950 10446 4002 10498
rect 19742 10446 19794 10498
rect 21870 10446 21922 10498
rect 22990 10446 23042 10498
rect 23326 10446 23378 10498
rect 27694 10446 27746 10498
rect 50878 10446 50930 10498
rect 7198 10334 7250 10386
rect 12238 10334 12290 10386
rect 32174 10334 32226 10386
rect 38446 10334 38498 10386
rect 38782 10334 38834 10386
rect 39454 10334 39506 10386
rect 45390 10334 45442 10386
rect 45614 10334 45666 10386
rect 45838 10334 45890 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 24446 9998 24498 10050
rect 2606 9886 2658 9938
rect 4734 9886 4786 9938
rect 8094 9886 8146 9938
rect 12238 9886 12290 9938
rect 16494 9886 16546 9938
rect 18622 9886 18674 9938
rect 19070 9886 19122 9938
rect 21982 9886 22034 9938
rect 32622 9886 32674 9938
rect 33070 9886 33122 9938
rect 38334 9886 38386 9938
rect 40462 9886 40514 9938
rect 41806 9886 41858 9938
rect 43934 9886 43986 9938
rect 45502 9886 45554 9938
rect 47630 9886 47682 9938
rect 52446 9886 52498 9938
rect 53454 9886 53506 9938
rect 55582 9886 55634 9938
rect 56814 9886 56866 9938
rect 1934 9774 1986 9826
rect 6974 9774 7026 9826
rect 7870 9774 7922 9826
rect 8542 9774 8594 9826
rect 9886 9774 9938 9826
rect 11006 9774 11058 9826
rect 12574 9774 12626 9826
rect 15710 9774 15762 9826
rect 22206 9774 22258 9826
rect 24670 9774 24722 9826
rect 24894 9774 24946 9826
rect 27470 9774 27522 9826
rect 27582 9774 27634 9826
rect 27806 9774 27858 9826
rect 29822 9774 29874 9826
rect 37662 9774 37714 9826
rect 41022 9774 41074 9826
rect 48302 9774 48354 9826
rect 49534 9774 49586 9826
rect 56366 9774 56418 9826
rect 6750 9662 6802 9714
rect 6862 9662 6914 9714
rect 8318 9662 8370 9714
rect 10782 9662 10834 9714
rect 11342 9662 11394 9714
rect 11902 9662 11954 9714
rect 27134 9662 27186 9714
rect 30494 9662 30546 9714
rect 50318 9662 50370 9714
rect 7422 9550 7474 9602
rect 9326 9550 9378 9602
rect 10222 9550 10274 9602
rect 11006 9550 11058 9602
rect 22542 9550 22594 9602
rect 24782 9550 24834 9602
rect 44382 9550 44434 9602
rect 48862 9550 48914 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 8206 9214 8258 9266
rect 10110 9214 10162 9266
rect 19070 9214 19122 9266
rect 26910 9214 26962 9266
rect 30718 9214 30770 9266
rect 45166 9214 45218 9266
rect 48078 9214 48130 9266
rect 5966 9102 6018 9154
rect 7646 9102 7698 9154
rect 8654 9102 8706 9154
rect 8878 9102 8930 9154
rect 9774 9102 9826 9154
rect 9998 9102 10050 9154
rect 13470 9102 13522 9154
rect 27470 9102 27522 9154
rect 27806 9102 27858 9154
rect 42590 9102 42642 9154
rect 48750 9102 48802 9154
rect 55358 9102 55410 9154
rect 4062 8990 4114 9042
rect 6190 8990 6242 9042
rect 7198 8990 7250 9042
rect 7422 8990 7474 9042
rect 7982 8990 8034 9042
rect 10558 8990 10610 9042
rect 12798 8990 12850 9042
rect 16046 8990 16098 9042
rect 20414 8990 20466 9042
rect 27134 8990 27186 9042
rect 39454 8990 39506 9042
rect 40238 8990 40290 9042
rect 40686 8990 40738 9042
rect 41806 8990 41858 9042
rect 50878 8990 50930 9042
rect 3278 8878 3330 8930
rect 3390 8878 3442 8930
rect 11006 8878 11058 8930
rect 15598 8878 15650 8930
rect 23214 8878 23266 8930
rect 27918 8878 27970 8930
rect 38670 8878 38722 8930
rect 39230 8878 39282 8930
rect 44718 8878 44770 8930
rect 51550 8878 51602 8930
rect 8990 8766 9042 8818
rect 10222 8766 10274 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 21758 8430 21810 8482
rect 22094 8430 22146 8482
rect 22878 8430 22930 8482
rect 27806 8430 27858 8482
rect 4958 8318 5010 8370
rect 6526 8318 6578 8370
rect 8654 8318 8706 8370
rect 16606 8318 16658 8370
rect 18734 8318 18786 8370
rect 24782 8318 24834 8370
rect 26910 8318 26962 8370
rect 28030 8318 28082 8370
rect 51886 8318 51938 8370
rect 52670 8318 52722 8370
rect 2158 8206 2210 8258
rect 5742 8206 5794 8258
rect 9662 8206 9714 8258
rect 10222 8206 10274 8258
rect 11006 8206 11058 8258
rect 11342 8206 11394 8258
rect 11566 8206 11618 8258
rect 11790 8206 11842 8258
rect 15822 8206 15874 8258
rect 20862 8206 20914 8258
rect 21870 8206 21922 8258
rect 22318 8206 22370 8258
rect 23998 8206 24050 8258
rect 44606 8206 44658 8258
rect 48974 8206 49026 8258
rect 49758 8206 49810 8258
rect 53566 8206 53618 8258
rect 53790 8206 53842 8258
rect 54014 8206 54066 8258
rect 54126 8206 54178 8258
rect 2830 8094 2882 8146
rect 10110 8094 10162 8146
rect 12014 8094 12066 8146
rect 42478 8094 42530 8146
rect 9214 7982 9266 8034
rect 9886 7982 9938 8034
rect 12126 7982 12178 8034
rect 19182 7982 19234 8034
rect 20638 7982 20690 8034
rect 20750 7982 20802 8034
rect 22990 7982 23042 8034
rect 23102 7982 23154 8034
rect 27470 7982 27522 8034
rect 38782 7982 38834 8034
rect 45502 7982 45554 8034
rect 47182 7982 47234 8034
rect 54126 7982 54178 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 2830 7646 2882 7698
rect 15934 7646 15986 7698
rect 30494 7646 30546 7698
rect 51774 7646 51826 7698
rect 55694 7646 55746 7698
rect 3166 7534 3218 7586
rect 3950 7534 4002 7586
rect 14702 7534 14754 7586
rect 22766 7534 22818 7586
rect 22990 7534 23042 7586
rect 24670 7534 24722 7586
rect 26238 7534 26290 7586
rect 43262 7534 43314 7586
rect 50430 7534 50482 7586
rect 54462 7534 54514 7586
rect 2606 7422 2658 7474
rect 2830 7422 2882 7474
rect 8990 7422 9042 7474
rect 10894 7422 10946 7474
rect 15486 7422 15538 7474
rect 19182 7422 19234 7474
rect 26574 7422 26626 7474
rect 29934 7422 29986 7474
rect 38222 7422 38274 7474
rect 39342 7422 39394 7474
rect 39790 7422 39842 7474
rect 42478 7422 42530 7474
rect 55246 7422 55298 7474
rect 10782 7310 10834 7362
rect 12574 7310 12626 7362
rect 19966 7310 20018 7362
rect 22094 7310 22146 7362
rect 22654 7310 22706 7362
rect 23662 7310 23714 7362
rect 24558 7310 24610 7362
rect 25566 7310 25618 7362
rect 27134 7310 27186 7362
rect 29262 7310 29314 7362
rect 38334 7310 38386 7362
rect 38558 7310 38610 7362
rect 39118 7310 39170 7362
rect 41918 7310 41970 7362
rect 45390 7310 45442 7362
rect 52334 7310 52386 7362
rect 10222 7198 10274 7250
rect 24446 7198 24498 7250
rect 26574 7198 26626 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 11902 6862 11954 6914
rect 27694 6862 27746 6914
rect 9214 6750 9266 6802
rect 11342 6750 11394 6802
rect 12238 6750 12290 6802
rect 22654 6750 22706 6802
rect 23886 6750 23938 6802
rect 26014 6750 26066 6802
rect 26798 6750 26850 6802
rect 38334 6750 38386 6802
rect 40462 6750 40514 6802
rect 49086 6750 49138 6802
rect 50430 6750 50482 6802
rect 52558 6750 52610 6802
rect 53342 6750 53394 6802
rect 2270 6638 2322 6690
rect 2718 6638 2770 6690
rect 4174 6638 4226 6690
rect 8542 6638 8594 6690
rect 12462 6638 12514 6690
rect 23214 6638 23266 6690
rect 27246 6638 27298 6690
rect 27470 6638 27522 6690
rect 27806 6638 27858 6690
rect 37662 6638 37714 6690
rect 46286 6638 46338 6690
rect 46958 6638 47010 6690
rect 49646 6638 49698 6690
rect 3726 6526 3778 6578
rect 2830 6414 2882 6466
rect 22094 6414 22146 6466
rect 40910 6414 40962 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 11790 6078 11842 6130
rect 22430 6078 22482 6130
rect 26238 6078 26290 6130
rect 40014 6078 40066 6130
rect 49422 6078 49474 6130
rect 52782 6078 52834 6130
rect 3950 5966 4002 6018
rect 11902 5966 11954 6018
rect 12126 5966 12178 6018
rect 19854 5966 19906 6018
rect 39230 5966 39282 6018
rect 39790 5966 39842 6018
rect 54126 5966 54178 6018
rect 4734 5854 4786 5906
rect 11454 5854 11506 5906
rect 19182 5854 19234 5906
rect 53342 5854 53394 5906
rect 1822 5742 1874 5794
rect 21982 5742 22034 5794
rect 56254 5742 56306 5794
rect 40126 5630 40178 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 41246 5182 41298 5234
rect 43374 5182 43426 5234
rect 55358 5182 55410 5234
rect 40574 5070 40626 5122
rect 43934 5070 43986 5122
rect 56142 5070 56194 5122
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 2494 3614 2546 3666
rect 22430 3614 22482 3666
rect 45614 3614 45666 3666
rect 1822 3502 1874 3554
rect 21982 3502 22034 3554
rect 44942 3502 44994 3554
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 5376 59200 5488 59800
rect 26880 59200 26992 59800
rect 49056 59200 49168 59800
rect 5404 56642 5460 59200
rect 5404 56590 5406 56642
rect 5458 56590 5460 56642
rect 5404 56578 5460 56590
rect 6412 56642 6468 56654
rect 6412 56590 6414 56642
rect 6466 56590 6468 56642
rect 5068 56084 5124 56094
rect 5740 56084 5796 56094
rect 5068 56082 5796 56084
rect 5068 56030 5070 56082
rect 5122 56030 5742 56082
rect 5794 56030 5796 56082
rect 5068 56028 5796 56030
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4172 51940 4228 51950
rect 2044 50708 2100 50718
rect 2044 50614 2100 50652
rect 4172 50706 4228 51884
rect 4956 51266 5012 51278
rect 4956 51214 4958 51266
rect 5010 51214 5012 51266
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4172 50654 4174 50706
rect 4226 50654 4228 50706
rect 4172 50642 4228 50654
rect 4284 50596 4340 50606
rect 4284 49810 4340 50540
rect 4956 50596 5012 51214
rect 5068 50708 5124 56028
rect 5740 56018 5796 56028
rect 6412 55970 6468 56590
rect 26908 56642 26964 59200
rect 26908 56590 26910 56642
rect 26962 56590 26964 56642
rect 26908 56578 26964 56590
rect 27804 56642 27860 56654
rect 27804 56590 27806 56642
rect 27858 56590 27860 56642
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 6412 55918 6414 55970
rect 6466 55918 6468 55970
rect 6412 55906 6468 55918
rect 27244 56082 27300 56094
rect 27244 56030 27246 56082
rect 27298 56030 27300 56082
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 8316 52164 8372 52174
rect 8316 52070 8372 52108
rect 8876 52164 8932 52174
rect 8428 51940 8484 51950
rect 8428 51846 8484 51884
rect 8540 51938 8596 51950
rect 8540 51886 8542 51938
rect 8594 51886 8596 51938
rect 8540 51828 8596 51886
rect 8540 51762 8596 51772
rect 5068 50642 5124 50652
rect 4956 50464 5012 50540
rect 6524 50596 6580 50606
rect 6524 50502 6580 50540
rect 7308 50482 7364 50494
rect 7308 50430 7310 50482
rect 7362 50430 7364 50482
rect 7308 50036 7364 50430
rect 7308 49970 7364 49980
rect 8652 50036 8708 50046
rect 8652 50034 8820 50036
rect 8652 49982 8654 50034
rect 8706 49982 8820 50034
rect 8652 49980 8820 49982
rect 8652 49970 8708 49980
rect 8764 49924 8820 49980
rect 8764 49858 8820 49868
rect 4284 49758 4286 49810
rect 4338 49758 4340 49810
rect 4284 49746 4340 49758
rect 8316 49810 8372 49822
rect 8652 49812 8708 49822
rect 8316 49758 8318 49810
rect 8370 49758 8372 49810
rect 4956 49698 5012 49710
rect 4956 49646 4958 49698
rect 5010 49646 5012 49698
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4956 48356 5012 49646
rect 7084 49698 7140 49710
rect 7084 49646 7086 49698
rect 7138 49646 7140 49698
rect 7084 49028 7140 49646
rect 7308 49028 7364 49038
rect 7084 48972 7308 49028
rect 7308 48934 7364 48972
rect 7532 49026 7588 49038
rect 7532 48974 7534 49026
rect 7586 48974 7588 49026
rect 7532 48692 7588 48974
rect 7532 48626 7588 48636
rect 7868 48802 7924 48814
rect 7868 48750 7870 48802
rect 7922 48750 7924 48802
rect 4956 48290 5012 48300
rect 7308 48356 7364 48366
rect 7308 48262 7364 48300
rect 7420 48244 7476 48254
rect 7420 48150 7476 48188
rect 7644 48244 7700 48254
rect 7868 48244 7924 48750
rect 7644 48242 7924 48244
rect 7644 48190 7646 48242
rect 7698 48190 7924 48242
rect 7644 48188 7924 48190
rect 7980 48804 8036 48814
rect 7644 48178 7700 48188
rect 7980 48132 8036 48748
rect 7756 48076 8036 48132
rect 8316 48692 8372 49758
rect 7756 48018 7812 48076
rect 7756 47966 7758 48018
rect 7810 47966 7812 48018
rect 7756 47954 7812 47966
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 7868 47572 7924 47582
rect 7644 47458 7700 47470
rect 7644 47406 7646 47458
rect 7698 47406 7700 47458
rect 7308 47234 7364 47246
rect 7308 47182 7310 47234
rect 7362 47182 7364 47234
rect 7308 47124 7364 47182
rect 7644 47236 7700 47406
rect 7644 47170 7700 47180
rect 7308 47058 7364 47068
rect 3500 46786 3556 46798
rect 3500 46734 3502 46786
rect 3554 46734 3556 46786
rect 2828 46004 2884 46014
rect 2828 45910 2884 45948
rect 3500 46004 3556 46734
rect 5740 46788 5796 46798
rect 5740 46694 5796 46732
rect 5068 46674 5124 46686
rect 5068 46622 5070 46674
rect 5122 46622 5124 46674
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 3500 45938 3556 45948
rect 4956 46004 5012 46014
rect 4956 45910 5012 45948
rect 2044 45892 2100 45902
rect 1932 45890 2100 45892
rect 1932 45838 2046 45890
rect 2098 45838 2100 45890
rect 1932 45836 2100 45838
rect 1932 44322 1988 45836
rect 2044 45826 2100 45836
rect 5068 45668 5124 46622
rect 7868 46562 7924 47516
rect 8316 47124 8372 48636
rect 8540 49810 8708 49812
rect 8540 49758 8654 49810
rect 8706 49758 8708 49810
rect 8540 49756 8708 49758
rect 8540 49028 8596 49756
rect 8652 49746 8708 49756
rect 8540 48802 8596 48972
rect 8764 48914 8820 48926
rect 8764 48862 8766 48914
rect 8818 48862 8820 48914
rect 8540 48750 8542 48802
rect 8594 48750 8596 48802
rect 8540 48580 8596 48750
rect 8652 48804 8708 48814
rect 8652 48710 8708 48748
rect 8764 48692 8820 48862
rect 8764 48626 8820 48636
rect 8876 48580 8932 52108
rect 9100 52164 9156 52174
rect 9100 52070 9156 52108
rect 19516 51940 19572 51950
rect 19292 51938 19572 51940
rect 19292 51886 19518 51938
rect 19570 51886 19572 51938
rect 19292 51884 19572 51886
rect 9324 51828 9380 51838
rect 8988 51380 9044 51390
rect 8988 51286 9044 51324
rect 9324 50708 9380 51772
rect 19292 51490 19348 51884
rect 19516 51874 19572 51884
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19292 51438 19294 51490
rect 19346 51438 19348 51490
rect 19292 51426 19348 51438
rect 9772 51380 9828 51390
rect 9772 51286 9828 51324
rect 14140 51380 14196 51390
rect 13244 51266 13300 51278
rect 13244 51214 13246 51266
rect 13298 51214 13300 51266
rect 9436 50708 9492 50718
rect 9324 50706 9492 50708
rect 9324 50654 9438 50706
rect 9490 50654 9492 50706
rect 9324 50652 9492 50654
rect 8988 49812 9044 49822
rect 9324 49812 9380 50652
rect 9436 50642 9492 50652
rect 12908 50706 12964 50718
rect 12908 50654 12910 50706
rect 12962 50654 12964 50706
rect 10108 50596 10164 50606
rect 10108 50502 10164 50540
rect 12012 50596 12068 50606
rect 10780 50482 10836 50494
rect 10780 50430 10782 50482
rect 10834 50430 10836 50482
rect 9884 50036 9940 50046
rect 9884 49942 9940 49980
rect 10780 50036 10836 50430
rect 10780 49970 10836 49980
rect 11676 50036 11732 50046
rect 11676 49942 11732 49980
rect 9772 49924 9828 49934
rect 9772 49830 9828 49868
rect 8988 49810 9380 49812
rect 8988 49758 8990 49810
rect 9042 49758 9380 49810
rect 8988 49756 9380 49758
rect 10108 49810 10164 49822
rect 10108 49758 10110 49810
rect 10162 49758 10164 49810
rect 8988 49746 9044 49756
rect 8540 48524 8708 48580
rect 8876 48524 9044 48580
rect 8652 48468 8708 48524
rect 8652 48412 8932 48468
rect 8540 48356 8596 48366
rect 8540 48354 8708 48356
rect 8540 48302 8542 48354
rect 8594 48302 8708 48354
rect 8540 48300 8708 48302
rect 8540 48290 8596 48300
rect 8540 48130 8596 48142
rect 8540 48078 8542 48130
rect 8594 48078 8596 48130
rect 8428 47346 8484 47358
rect 8428 47294 8430 47346
rect 8482 47294 8484 47346
rect 8428 47236 8484 47294
rect 8428 47170 8484 47180
rect 8316 47058 8372 47068
rect 8540 46674 8596 48078
rect 8652 47572 8708 48300
rect 8652 47458 8708 47516
rect 8652 47406 8654 47458
rect 8706 47406 8708 47458
rect 8652 47394 8708 47406
rect 8764 48018 8820 48030
rect 8764 47966 8766 48018
rect 8818 47966 8820 48018
rect 8764 47236 8820 47966
rect 8876 47458 8932 48412
rect 8876 47406 8878 47458
rect 8930 47406 8932 47458
rect 8876 47394 8932 47406
rect 8988 48244 9044 48524
rect 8988 47236 9044 48188
rect 9100 47458 9156 49756
rect 10108 49588 10164 49758
rect 11900 49812 11956 49822
rect 11900 49718 11956 49756
rect 9660 48244 9716 48254
rect 9660 48150 9716 48188
rect 9100 47406 9102 47458
rect 9154 47406 9156 47458
rect 9100 47394 9156 47406
rect 10108 47346 10164 49532
rect 11564 49588 11620 49598
rect 11564 49494 11620 49532
rect 10780 48132 10836 48142
rect 10108 47294 10110 47346
rect 10162 47294 10164 47346
rect 10108 47282 10164 47294
rect 10444 47348 10500 47358
rect 10444 47346 10724 47348
rect 10444 47294 10446 47346
rect 10498 47294 10724 47346
rect 10444 47292 10724 47294
rect 10444 47282 10500 47292
rect 8764 47170 8820 47180
rect 8876 47180 9044 47236
rect 9212 47236 9268 47246
rect 10220 47236 10276 47246
rect 9212 47234 9828 47236
rect 9212 47182 9214 47234
rect 9266 47182 9828 47234
rect 9212 47180 9828 47182
rect 8540 46622 8542 46674
rect 8594 46622 8596 46674
rect 8540 46610 8596 46622
rect 8652 47012 8708 47022
rect 8652 46674 8708 46956
rect 8652 46622 8654 46674
rect 8706 46622 8708 46674
rect 8652 46610 8708 46622
rect 8876 46674 8932 47180
rect 9212 47170 9268 47180
rect 8988 46788 9044 46798
rect 8988 46694 9044 46732
rect 8876 46622 8878 46674
rect 8930 46622 8932 46674
rect 7868 46510 7870 46562
rect 7922 46510 7924 46562
rect 7868 46498 7924 46510
rect 8876 46452 8932 46622
rect 8876 46396 9268 46452
rect 4956 45332 5012 45342
rect 5068 45332 5124 45612
rect 4956 45330 5124 45332
rect 4956 45278 4958 45330
rect 5010 45278 5124 45330
rect 4956 45276 5124 45278
rect 5404 46004 5460 46014
rect 4956 45266 5012 45276
rect 2716 45218 2772 45230
rect 2716 45166 2718 45218
rect 2770 45166 2772 45218
rect 2604 44436 2660 44446
rect 2716 44436 2772 45166
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 2604 44434 2772 44436
rect 2604 44382 2606 44434
rect 2658 44382 2772 44434
rect 2604 44380 2772 44382
rect 4732 44434 4788 44446
rect 4732 44382 4734 44434
rect 4786 44382 4788 44434
rect 2604 44370 2660 44380
rect 1932 44270 1934 44322
rect 1986 44270 1988 44322
rect 1932 42756 1988 44270
rect 4172 43764 4228 43774
rect 2828 43650 2884 43662
rect 2828 43598 2830 43650
rect 2882 43598 2884 43650
rect 2828 42866 2884 43598
rect 2828 42814 2830 42866
rect 2882 42814 2884 42866
rect 2828 42802 2884 42814
rect 2156 42756 2212 42766
rect 1932 42754 2212 42756
rect 1932 42702 2158 42754
rect 2210 42702 2212 42754
rect 1932 42700 2212 42702
rect 2156 41972 2212 42700
rect 1932 41916 2156 41972
rect 1932 41186 1988 41916
rect 2156 41906 2212 41916
rect 2716 42082 2772 42094
rect 2716 42030 2718 42082
rect 2770 42030 2772 42082
rect 2604 41300 2660 41310
rect 2716 41300 2772 42030
rect 2604 41298 2772 41300
rect 2604 41246 2606 41298
rect 2658 41246 2772 41298
rect 2604 41244 2772 41246
rect 2604 41234 2660 41244
rect 1932 41134 1934 41186
rect 1986 41134 1988 41186
rect 1932 41122 1988 41134
rect 3052 30884 3108 30894
rect 3052 30790 3108 30828
rect 4172 28756 4228 43708
rect 4732 43708 4788 44382
rect 4732 43652 5236 43708
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4956 42866 5012 42878
rect 4956 42814 4958 42866
rect 5010 42814 5012 42866
rect 4956 42084 5012 42814
rect 4956 42028 5124 42084
rect 4396 41972 4452 41982
rect 4396 41878 4452 41916
rect 4956 41860 5012 41870
rect 4844 41858 5012 41860
rect 4844 41806 4958 41858
rect 5010 41806 5012 41858
rect 4844 41804 5012 41806
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4732 41300 4788 41310
rect 4844 41300 4900 41804
rect 4956 41794 5012 41804
rect 5068 41860 5124 42028
rect 5180 41970 5236 43652
rect 5180 41918 5182 41970
rect 5234 41918 5236 41970
rect 5180 41906 5236 41918
rect 5404 41970 5460 45948
rect 9212 46004 9268 46396
rect 9212 46002 9716 46004
rect 9212 45950 9214 46002
rect 9266 45950 9716 46002
rect 9212 45948 9716 45950
rect 9212 45938 9268 45948
rect 5628 45668 5684 45678
rect 5628 45574 5684 45612
rect 5852 45668 5908 45678
rect 5404 41918 5406 41970
rect 5458 41918 5460 41970
rect 5404 41906 5460 41918
rect 5852 44434 5908 45612
rect 8092 45668 8148 45678
rect 8092 45574 8148 45612
rect 7308 45218 7364 45230
rect 7308 45166 7310 45218
rect 7362 45166 7364 45218
rect 5852 44382 5854 44434
rect 5906 44382 5908 44434
rect 5852 44324 5908 44382
rect 7196 44436 7252 44446
rect 7308 44436 7364 45166
rect 9660 44548 9716 45948
rect 9772 45218 9828 47180
rect 9884 46676 9940 46686
rect 9884 46582 9940 46620
rect 10220 45892 10276 47180
rect 10556 46562 10612 46574
rect 10556 46510 10558 46562
rect 10610 46510 10612 46562
rect 10332 46116 10388 46126
rect 10556 46116 10612 46510
rect 10332 46114 10612 46116
rect 10332 46062 10334 46114
rect 10386 46062 10612 46114
rect 10332 46060 10612 46062
rect 10332 46050 10388 46060
rect 10444 45892 10500 45902
rect 10668 45892 10724 47292
rect 10780 46114 10836 48076
rect 11900 47236 11956 47246
rect 11900 47142 11956 47180
rect 12012 46676 12068 50540
rect 12460 50036 12516 50046
rect 12460 49922 12516 49980
rect 12460 49870 12462 49922
rect 12514 49870 12516 49922
rect 12460 49252 12516 49870
rect 12684 49924 12740 49934
rect 12908 49924 12964 50654
rect 13244 50596 13300 51214
rect 13244 50530 13300 50540
rect 13692 50706 13748 50718
rect 13692 50654 13694 50706
rect 13746 50654 13748 50706
rect 13692 50036 13748 50654
rect 13692 49970 13748 49980
rect 13916 50484 13972 50494
rect 12684 49922 12964 49924
rect 12684 49870 12686 49922
rect 12738 49870 12964 49922
rect 12684 49868 12964 49870
rect 13916 49922 13972 50428
rect 13916 49870 13918 49922
rect 13970 49870 13972 49922
rect 12684 49812 12740 49868
rect 13916 49858 13972 49870
rect 12572 49252 12628 49262
rect 12236 49250 12628 49252
rect 12236 49198 12574 49250
rect 12626 49198 12628 49250
rect 12236 49196 12628 49198
rect 12236 47458 12292 49196
rect 12572 49186 12628 49196
rect 12348 49026 12404 49038
rect 12348 48974 12350 49026
rect 12402 48974 12404 49026
rect 12348 48804 12404 48974
rect 12684 48804 12740 49756
rect 13356 49810 13412 49822
rect 13356 49758 13358 49810
rect 13410 49758 13412 49810
rect 12796 49700 12852 49710
rect 13356 49700 13412 49758
rect 12796 49698 13412 49700
rect 12796 49646 12798 49698
rect 12850 49646 13412 49698
rect 12796 49644 13412 49646
rect 12796 49634 12852 49644
rect 13580 49588 13636 49598
rect 12348 48748 12740 48804
rect 12236 47406 12238 47458
rect 12290 47406 12292 47458
rect 12236 47394 12292 47406
rect 12460 48244 12516 48254
rect 12460 47346 12516 48188
rect 12572 48242 12628 48254
rect 12572 48190 12574 48242
rect 12626 48190 12628 48242
rect 12572 47572 12628 48190
rect 12684 48020 12740 48748
rect 12908 48804 12964 48814
rect 12908 48710 12964 48748
rect 13132 48804 13188 48814
rect 12796 48244 12852 48254
rect 12796 48150 12852 48188
rect 13132 48242 13188 48748
rect 13580 48356 13636 49532
rect 13804 49586 13860 49598
rect 13804 49534 13806 49586
rect 13858 49534 13860 49586
rect 13804 48804 13860 49534
rect 13804 48738 13860 48748
rect 14028 48804 14084 48814
rect 13580 48300 13860 48356
rect 13132 48190 13134 48242
rect 13186 48190 13188 48242
rect 13132 48178 13188 48190
rect 13244 48244 13300 48254
rect 12908 48132 12964 48142
rect 12908 48038 12964 48076
rect 12684 47964 12852 48020
rect 12572 47516 12740 47572
rect 12460 47294 12462 47346
rect 12514 47294 12516 47346
rect 12460 47282 12516 47294
rect 12684 47458 12740 47516
rect 12684 47406 12686 47458
rect 12738 47406 12740 47458
rect 12012 46610 12068 46620
rect 12684 46562 12740 47406
rect 12796 47458 12852 47964
rect 12796 47406 12798 47458
rect 12850 47406 12852 47458
rect 12796 47394 12852 47406
rect 12684 46510 12686 46562
rect 12738 46510 12740 46562
rect 12684 46498 12740 46510
rect 12908 46676 12964 46686
rect 10780 46062 10782 46114
rect 10834 46062 10836 46114
rect 10780 46050 10836 46062
rect 10220 45890 10500 45892
rect 10220 45838 10446 45890
rect 10498 45838 10500 45890
rect 10220 45836 10500 45838
rect 10444 45826 10500 45836
rect 10556 45890 10724 45892
rect 10556 45838 10670 45890
rect 10722 45838 10724 45890
rect 10556 45836 10724 45838
rect 10556 45330 10612 45836
rect 10668 45826 10724 45836
rect 12908 46002 12964 46620
rect 13244 46562 13300 48188
rect 13244 46510 13246 46562
rect 13298 46510 13300 46562
rect 13244 46498 13300 46510
rect 13692 46564 13748 46574
rect 12908 45950 12910 46002
rect 12962 45950 12964 46002
rect 12908 45892 12964 45950
rect 13580 46004 13636 46014
rect 13580 45910 13636 45948
rect 12908 45826 12964 45836
rect 10556 45278 10558 45330
rect 10610 45278 10612 45330
rect 10556 45266 10612 45278
rect 9772 45166 9774 45218
rect 9826 45166 9828 45218
rect 9772 45154 9828 45166
rect 9884 45108 9940 45118
rect 9772 44548 9828 44558
rect 9660 44546 9828 44548
rect 9660 44494 9774 44546
rect 9826 44494 9828 44546
rect 9660 44492 9828 44494
rect 9772 44482 9828 44492
rect 7196 44434 7364 44436
rect 7196 44382 7198 44434
rect 7250 44382 7364 44434
rect 7196 44380 7364 44382
rect 9324 44434 9380 44446
rect 9324 44382 9326 44434
rect 9378 44382 9380 44434
rect 7196 44370 7252 44380
rect 5852 43650 5908 44268
rect 6412 44324 6468 44334
rect 6412 44230 6468 44268
rect 5852 43598 5854 43650
rect 5906 43598 5908 43650
rect 5852 41972 5908 43598
rect 8316 43538 8372 43550
rect 8316 43486 8318 43538
rect 8370 43486 8372 43538
rect 8316 43428 8372 43486
rect 9324 43540 9380 44382
rect 9884 44210 9940 45052
rect 9996 45106 10052 45118
rect 9996 45054 9998 45106
rect 10050 45054 10052 45106
rect 9996 44324 10052 45054
rect 10220 45106 10276 45118
rect 10220 45054 10222 45106
rect 10274 45054 10276 45106
rect 9996 44258 10052 44268
rect 10108 44324 10164 44334
rect 10220 44324 10276 45054
rect 10444 45108 10500 45118
rect 10444 45014 10500 45052
rect 13692 44994 13748 46508
rect 13804 45330 13860 48300
rect 13916 48244 13972 48254
rect 13916 48150 13972 48188
rect 14028 48130 14084 48748
rect 14028 48078 14030 48130
rect 14082 48078 14084 48130
rect 14028 48066 14084 48078
rect 14140 47458 14196 51324
rect 18508 51378 18564 51390
rect 18508 51326 18510 51378
rect 18562 51326 18564 51378
rect 14364 50596 14420 50606
rect 14364 49026 14420 50540
rect 16604 50594 16660 50606
rect 16604 50542 16606 50594
rect 16658 50542 16660 50594
rect 15820 50484 15876 50494
rect 15820 50390 15876 50428
rect 16604 50484 16660 50542
rect 16604 50418 16660 50428
rect 17052 50484 17108 50494
rect 17052 50390 17108 50428
rect 17948 50484 18004 50494
rect 16380 49924 16436 49934
rect 15148 49922 16436 49924
rect 15148 49870 16382 49922
rect 16434 49870 16436 49922
rect 15148 49868 16436 49870
rect 15148 49138 15204 49868
rect 16380 49858 16436 49868
rect 15148 49086 15150 49138
rect 15202 49086 15204 49138
rect 15148 49074 15204 49086
rect 17276 49138 17332 49150
rect 17276 49086 17278 49138
rect 17330 49086 17332 49138
rect 14364 48974 14366 49026
rect 14418 48974 14420 49026
rect 14364 48962 14420 48974
rect 17276 49028 17332 49086
rect 17276 48962 17332 48972
rect 17948 49028 18004 50428
rect 18508 50484 18564 51326
rect 21420 51268 21476 51278
rect 21980 51268 22036 51278
rect 21420 51266 21812 51268
rect 21420 51214 21422 51266
rect 21474 51214 21812 51266
rect 21420 51212 21812 51214
rect 21420 51202 21476 51212
rect 18508 50418 18564 50428
rect 19628 50484 19684 50494
rect 19628 49812 19684 50428
rect 21644 50372 21700 50382
rect 20748 50370 21700 50372
rect 20748 50318 21646 50370
rect 21698 50318 21700 50370
rect 20748 50316 21700 50318
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19964 49924 20020 49934
rect 19964 49812 20020 49868
rect 20748 49922 20804 50316
rect 21644 50306 21700 50316
rect 20748 49870 20750 49922
rect 20802 49870 20804 49922
rect 20748 49858 20804 49870
rect 20972 49924 21028 49934
rect 19628 49810 20020 49812
rect 19628 49758 19966 49810
rect 20018 49758 20020 49810
rect 19628 49756 20020 49758
rect 19964 49746 20020 49756
rect 20748 49140 20804 49150
rect 20748 49046 20804 49084
rect 17948 49026 18116 49028
rect 17948 48974 17950 49026
rect 18002 48974 18116 49026
rect 17948 48972 18116 48974
rect 17948 48962 18004 48972
rect 17612 48130 17668 48142
rect 17612 48078 17614 48130
rect 17666 48078 17668 48130
rect 14140 47406 14142 47458
rect 14194 47406 14196 47458
rect 14140 46788 14196 47406
rect 14140 46004 14196 46732
rect 14140 45938 14196 45948
rect 14252 48018 14308 48030
rect 14252 47966 14254 48018
rect 14306 47966 14308 48018
rect 13804 45278 13806 45330
rect 13858 45278 13860 45330
rect 13804 45266 13860 45278
rect 13916 45892 13972 45902
rect 13692 44942 13694 44994
rect 13746 44942 13748 44994
rect 13692 44930 13748 44942
rect 10108 44322 10276 44324
rect 10108 44270 10110 44322
rect 10162 44270 10276 44322
rect 10108 44268 10276 44270
rect 10332 44324 10388 44334
rect 9884 44158 9886 44210
rect 9938 44158 9940 44210
rect 9884 43762 9940 44158
rect 9884 43710 9886 43762
rect 9938 43710 9940 43762
rect 9884 43698 9940 43710
rect 9324 43474 9380 43484
rect 8316 43362 8372 43372
rect 6188 43316 6244 43326
rect 5068 41794 5124 41804
rect 5628 41860 5684 41870
rect 5628 41766 5684 41804
rect 4732 41298 4900 41300
rect 4732 41246 4734 41298
rect 4786 41246 4900 41298
rect 4732 41244 4900 41246
rect 5740 41300 5796 41310
rect 5852 41300 5908 41916
rect 6076 42754 6132 42766
rect 6076 42702 6078 42754
rect 6130 42702 6132 42754
rect 6076 41972 6132 42702
rect 6076 41906 6132 41916
rect 6076 41748 6132 41758
rect 6188 41748 6244 43260
rect 9884 43316 9940 43326
rect 9884 43222 9940 43260
rect 9996 43314 10052 43326
rect 9996 43262 9998 43314
rect 10050 43262 10052 43314
rect 9100 42980 9156 42990
rect 8876 42978 9156 42980
rect 8876 42926 9102 42978
rect 9154 42926 9156 42978
rect 8876 42924 9156 42926
rect 8876 42866 8932 42924
rect 9100 42914 9156 42924
rect 9772 42980 9828 42990
rect 9996 42980 10052 43262
rect 9772 42978 10052 42980
rect 9772 42926 9774 42978
rect 9826 42926 10052 42978
rect 9772 42924 10052 42926
rect 10108 42980 10164 44268
rect 10332 43708 10388 44268
rect 13804 44324 13860 44334
rect 13916 44324 13972 45836
rect 14028 45220 14084 45230
rect 14252 45220 14308 47966
rect 16828 47346 16884 47358
rect 16828 47294 16830 47346
rect 16882 47294 16884 47346
rect 16828 46900 16884 47294
rect 15036 46788 15092 46798
rect 14476 45892 14532 45902
rect 14476 45798 14532 45836
rect 14028 45218 14308 45220
rect 14028 45166 14030 45218
rect 14082 45166 14308 45218
rect 14028 45164 14308 45166
rect 14028 45154 14084 45164
rect 13804 44322 13972 44324
rect 13804 44270 13806 44322
rect 13858 44270 13972 44322
rect 13804 44268 13972 44270
rect 13804 44258 13860 44268
rect 14476 44212 14532 44222
rect 13916 44210 14532 44212
rect 13916 44158 14478 44210
rect 14530 44158 14532 44210
rect 13916 44156 14532 44158
rect 13804 43764 13860 43774
rect 13916 43764 13972 44156
rect 14476 44146 14532 44156
rect 13804 43762 13972 43764
rect 13804 43710 13806 43762
rect 13858 43710 13972 43762
rect 13804 43708 13972 43710
rect 10332 43652 10500 43708
rect 13804 43698 13860 43708
rect 10220 43540 10276 43550
rect 10220 43446 10276 43484
rect 9772 42914 9828 42924
rect 10108 42914 10164 42924
rect 8876 42814 8878 42866
rect 8930 42814 8932 42866
rect 8876 42802 8932 42814
rect 9996 42754 10052 42766
rect 9996 42702 9998 42754
rect 10050 42702 10052 42754
rect 6748 42642 6804 42654
rect 6748 42590 6750 42642
rect 6802 42590 6804 42642
rect 6748 42196 6804 42590
rect 9324 42530 9380 42542
rect 9324 42478 9326 42530
rect 9378 42478 9380 42530
rect 6860 42196 6916 42206
rect 6748 42194 6916 42196
rect 6748 42142 6862 42194
rect 6914 42142 6916 42194
rect 6748 42140 6916 42142
rect 6860 42130 6916 42140
rect 6076 41746 6244 41748
rect 6076 41694 6078 41746
rect 6130 41694 6244 41746
rect 6076 41692 6244 41694
rect 8428 41972 8484 41982
rect 6076 41682 6132 41692
rect 5740 41298 5908 41300
rect 5740 41246 5742 41298
rect 5794 41246 5908 41298
rect 5740 41244 5908 41246
rect 4732 41234 4788 41244
rect 5740 41234 5796 41244
rect 8428 41186 8484 41916
rect 9324 41972 9380 42478
rect 9324 41906 9380 41916
rect 9996 41972 10052 42702
rect 9996 41906 10052 41916
rect 10332 41972 10388 41982
rect 10332 41858 10388 41916
rect 10332 41806 10334 41858
rect 10386 41806 10388 41858
rect 10332 41794 10388 41806
rect 10444 41300 10500 43652
rect 10780 43428 10836 43438
rect 10780 43334 10836 43372
rect 15036 43428 15092 46732
rect 16156 46674 16212 46686
rect 16156 46622 16158 46674
rect 16210 46622 16212 46674
rect 15372 46564 15428 46574
rect 15372 46470 15428 46508
rect 15260 45778 15316 45790
rect 15260 45726 15262 45778
rect 15314 45726 15316 45778
rect 15260 45332 15316 45726
rect 16156 45444 16212 46622
rect 16828 45892 16884 46844
rect 17612 46900 17668 48078
rect 17612 46806 17668 46844
rect 16940 46788 16996 46798
rect 16940 46694 16996 46732
rect 17388 46116 17444 46126
rect 17388 46002 17444 46060
rect 17388 45950 17390 46002
rect 17442 45950 17444 46002
rect 17388 45938 17444 45950
rect 16828 45826 16884 45836
rect 17164 45892 17220 45902
rect 16380 45444 16436 45454
rect 16156 45388 16380 45444
rect 15260 45266 15316 45276
rect 16380 45330 16436 45388
rect 16380 45278 16382 45330
rect 16434 45278 16436 45330
rect 16380 45266 16436 45278
rect 16604 44434 16660 44446
rect 16604 44382 16606 44434
rect 16658 44382 16660 44434
rect 16604 43708 16660 44382
rect 17164 44434 17220 45836
rect 18060 45890 18116 48972
rect 18620 48914 18676 48926
rect 18620 48862 18622 48914
rect 18674 48862 18676 48914
rect 18620 48468 18676 48862
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 18732 48468 18788 48478
rect 18620 48466 18788 48468
rect 18620 48414 18734 48466
rect 18786 48414 18788 48466
rect 18620 48412 18788 48414
rect 18732 48402 18788 48412
rect 20972 48466 21028 49868
rect 21756 49700 21812 51212
rect 21980 51266 23380 51268
rect 21980 51214 21982 51266
rect 22034 51214 23380 51266
rect 21980 51212 23380 51214
rect 21980 49924 22036 51212
rect 23324 50034 23380 51212
rect 26236 51266 26292 51278
rect 26236 51214 26238 51266
rect 26290 51214 26292 51266
rect 24444 50594 24500 50606
rect 24444 50542 24446 50594
rect 24498 50542 24500 50594
rect 24444 50484 24500 50542
rect 24444 50418 24500 50428
rect 25116 50482 25172 50494
rect 25116 50430 25118 50482
rect 25170 50430 25172 50482
rect 23324 49982 23326 50034
rect 23378 49982 23380 50034
rect 23324 49970 23380 49982
rect 21980 49858 22036 49868
rect 24892 49924 24948 49934
rect 22876 49700 22932 49710
rect 21756 49644 22148 49700
rect 22092 49250 22148 49644
rect 22092 49198 22094 49250
rect 22146 49198 22148 49250
rect 22092 49186 22148 49198
rect 22316 49698 22932 49700
rect 22316 49646 22878 49698
rect 22930 49646 22932 49698
rect 22316 49644 22932 49646
rect 22316 49250 22372 49644
rect 22876 49634 22932 49644
rect 24892 49698 24948 49868
rect 24892 49646 24894 49698
rect 24946 49646 24948 49698
rect 22316 49198 22318 49250
rect 22370 49198 22372 49250
rect 22316 49186 22372 49198
rect 24220 49588 24276 49598
rect 21868 49140 21924 49150
rect 21868 49046 21924 49084
rect 22988 49140 23044 49150
rect 22988 49046 23044 49084
rect 21644 49028 21700 49038
rect 21644 48934 21700 48972
rect 20972 48414 20974 48466
rect 21026 48414 21028 48466
rect 20972 48402 21028 48414
rect 22204 48802 22260 48814
rect 22204 48750 22206 48802
rect 22258 48750 22260 48802
rect 21644 47684 21700 47694
rect 21644 47590 21700 47628
rect 22204 47570 22260 48750
rect 22204 47518 22206 47570
rect 22258 47518 22260 47570
rect 22204 47506 22260 47518
rect 23212 48356 23268 48366
rect 23212 47684 23268 48300
rect 21980 47458 22036 47470
rect 21980 47406 21982 47458
rect 22034 47406 22036 47458
rect 19516 47236 19572 47246
rect 18732 47234 19572 47236
rect 18732 47182 19518 47234
rect 19570 47182 19572 47234
rect 18732 47180 19572 47182
rect 18396 46788 18452 46798
rect 18396 46674 18452 46732
rect 18396 46622 18398 46674
rect 18450 46622 18452 46674
rect 18396 46610 18452 46622
rect 18732 46002 18788 47180
rect 19516 47170 19572 47180
rect 20748 47234 20804 47246
rect 20748 47182 20750 47234
rect 20802 47182 20804 47234
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 18732 45950 18734 46002
rect 18786 45950 18788 46002
rect 18732 45938 18788 45950
rect 18060 45838 18062 45890
rect 18114 45838 18116 45890
rect 18060 45444 18116 45838
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20188 45444 20244 45454
rect 17724 45332 17780 45342
rect 17724 45238 17780 45276
rect 17164 44382 17166 44434
rect 17218 44382 17220 44434
rect 17164 44370 17220 44382
rect 15708 43652 16660 43708
rect 15260 43540 15316 43550
rect 14252 42980 14308 42990
rect 14252 42886 14308 42924
rect 14588 42980 14644 42990
rect 14588 42886 14644 42924
rect 12908 42868 12964 42878
rect 12908 42774 12964 42812
rect 14812 42756 14868 42766
rect 14812 42662 14868 42700
rect 8428 41134 8430 41186
rect 8482 41134 8484 41186
rect 8428 41122 8484 41134
rect 10332 41244 10500 41300
rect 10780 42642 10836 42654
rect 10780 42590 10782 42642
rect 10834 42590 10836 42642
rect 9100 41076 9156 41086
rect 9100 41074 9828 41076
rect 9100 41022 9102 41074
rect 9154 41022 9828 41074
rect 9100 41020 9828 41022
rect 9100 41010 9156 41020
rect 9772 40626 9828 41020
rect 9772 40574 9774 40626
rect 9826 40574 9828 40626
rect 9772 40562 9828 40574
rect 5852 40516 5908 40526
rect 5628 40514 5908 40516
rect 5628 40462 5854 40514
rect 5906 40462 5908 40514
rect 5628 40460 5908 40462
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 5628 38946 5684 40460
rect 5852 40450 5908 40460
rect 8092 40290 8148 40302
rect 8092 40238 8094 40290
rect 8146 40238 8148 40290
rect 5628 38894 5630 38946
rect 5682 38894 5684 38946
rect 5628 38882 5684 38894
rect 7644 39620 7700 39630
rect 8092 39620 8148 40238
rect 7644 39618 8148 39620
rect 7644 39566 7646 39618
rect 7698 39566 8148 39618
rect 7644 39564 8148 39566
rect 4956 38834 5012 38846
rect 4956 38782 4958 38834
rect 5010 38782 5012 38834
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4956 37268 5012 38782
rect 7644 37492 7700 39564
rect 8316 39508 8372 39518
rect 8316 39506 8596 39508
rect 8316 39454 8318 39506
rect 8370 39454 8596 39506
rect 8316 39452 8596 39454
rect 8316 39442 8372 39452
rect 8540 39058 8596 39452
rect 8540 39006 8542 39058
rect 8594 39006 8596 39058
rect 8540 38994 8596 39006
rect 10332 39058 10388 41244
rect 10780 41076 10836 42590
rect 13580 42530 13636 42542
rect 13580 42478 13582 42530
rect 13634 42478 13636 42530
rect 11676 41972 11732 41982
rect 11228 41300 11284 41310
rect 11228 41298 11396 41300
rect 11228 41246 11230 41298
rect 11282 41246 11396 41298
rect 11228 41244 11396 41246
rect 11228 41234 11284 41244
rect 10780 41010 10836 41020
rect 10444 39730 10500 39742
rect 10444 39678 10446 39730
rect 10498 39678 10500 39730
rect 10444 39172 10500 39678
rect 10892 39394 10948 39406
rect 10892 39342 10894 39394
rect 10946 39342 10948 39394
rect 10444 39116 10836 39172
rect 10332 39006 10334 39058
rect 10386 39006 10388 39058
rect 10332 38994 10388 39006
rect 9884 38946 9940 38958
rect 9884 38894 9886 38946
rect 9938 38894 9940 38946
rect 7756 38836 7812 38846
rect 7756 38722 7812 38780
rect 9772 38836 9828 38846
rect 9772 38742 9828 38780
rect 7756 38670 7758 38722
rect 7810 38670 7812 38722
rect 7756 38658 7812 38670
rect 9884 38164 9940 38894
rect 10780 38834 10836 39116
rect 10780 38782 10782 38834
rect 10834 38782 10836 38834
rect 10780 38770 10836 38782
rect 8652 38108 9940 38164
rect 8316 38052 8372 38062
rect 8316 37958 8372 37996
rect 7868 37492 7924 37502
rect 7644 37436 7868 37492
rect 5404 37268 5460 37278
rect 4956 37266 5460 37268
rect 4956 37214 5406 37266
rect 5458 37214 5460 37266
rect 4956 37212 5460 37214
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4508 35700 4564 35710
rect 4508 35606 4564 35644
rect 5404 35700 5460 37212
rect 6188 37156 6244 37166
rect 6188 37154 6468 37156
rect 6188 37102 6190 37154
rect 6242 37102 6468 37154
rect 6188 37100 6468 37102
rect 6188 37090 6244 37100
rect 6412 36370 6468 37100
rect 7756 36708 7812 36718
rect 7756 36614 7812 36652
rect 7532 36372 7588 36382
rect 6412 36318 6414 36370
rect 6466 36318 6468 36370
rect 6412 36306 6468 36318
rect 7308 36370 7588 36372
rect 7308 36318 7534 36370
rect 7586 36318 7588 36370
rect 7308 36316 7588 36318
rect 5404 35634 5460 35644
rect 5740 36258 5796 36270
rect 5740 36206 5742 36258
rect 5794 36206 5796 36258
rect 5180 35586 5236 35598
rect 5180 35534 5182 35586
rect 5234 35534 5236 35586
rect 5180 35476 5236 35534
rect 5740 35476 5796 36206
rect 7308 35586 7364 36316
rect 7532 36306 7588 36316
rect 7756 35700 7812 35710
rect 7868 35700 7924 37436
rect 8316 37154 8372 37166
rect 8316 37102 8318 37154
rect 8370 37102 8372 37154
rect 8316 36708 8372 37102
rect 8316 36642 8372 36652
rect 8652 36706 8708 38108
rect 8988 37938 9044 37950
rect 8988 37886 8990 37938
rect 9042 37886 9044 37938
rect 8764 37492 8820 37502
rect 8988 37492 9044 37886
rect 8820 37436 9044 37492
rect 10892 37492 10948 39342
rect 11340 38946 11396 41244
rect 11676 41188 11732 41916
rect 13580 41972 13636 42478
rect 13580 41906 13636 41916
rect 15036 41972 15092 43372
rect 11676 40626 11732 41132
rect 12348 41188 12404 41198
rect 11788 41076 11844 41086
rect 11788 40982 11844 41020
rect 11676 40574 11678 40626
rect 11730 40574 11732 40626
rect 11676 40562 11732 40574
rect 12348 40402 12404 41132
rect 13692 40962 13748 40974
rect 13692 40910 13694 40962
rect 13746 40910 13748 40962
rect 13020 40516 13076 40526
rect 13020 40422 13076 40460
rect 13692 40516 13748 40910
rect 13692 40450 13748 40460
rect 12348 40350 12350 40402
rect 12402 40350 12404 40402
rect 12348 39732 12404 40350
rect 15036 40404 15092 41916
rect 12460 39732 12516 39742
rect 12348 39730 12852 39732
rect 12348 39678 12462 39730
rect 12514 39678 12852 39730
rect 12348 39676 12852 39678
rect 12460 39666 12516 39676
rect 11340 38894 11342 38946
rect 11394 38894 11396 38946
rect 11340 38882 11396 38894
rect 12236 38948 12292 38958
rect 12236 38946 12628 38948
rect 12236 38894 12238 38946
rect 12290 38894 12628 38946
rect 12236 38892 12628 38894
rect 12236 38882 12292 38892
rect 8764 37398 8820 37436
rect 10892 37426 10948 37436
rect 11228 37492 11284 37502
rect 11228 37398 11284 37436
rect 11788 37492 11844 37502
rect 10108 37380 10164 37390
rect 10108 37378 10836 37380
rect 10108 37326 10110 37378
rect 10162 37326 10836 37378
rect 10108 37324 10836 37326
rect 10108 37314 10164 37324
rect 10780 36932 10836 37324
rect 11788 37266 11844 37436
rect 12572 37378 12628 38892
rect 12796 38834 12852 39676
rect 13804 39396 13860 39406
rect 13580 39394 13860 39396
rect 13580 39342 13806 39394
rect 13858 39342 13860 39394
rect 13580 39340 13860 39342
rect 13580 38946 13636 39340
rect 13804 39330 13860 39340
rect 13580 38894 13582 38946
rect 13634 38894 13636 38946
rect 13580 38882 13636 38894
rect 12796 38782 12798 38834
rect 12850 38782 12852 38834
rect 12796 38770 12852 38782
rect 12684 38164 12740 38174
rect 12684 38070 12740 38108
rect 13356 38164 13412 38174
rect 12572 37326 12574 37378
rect 12626 37326 12628 37378
rect 12572 37314 12628 37326
rect 11788 37214 11790 37266
rect 11842 37214 11844 37266
rect 11788 37202 11844 37214
rect 10780 36876 11284 36932
rect 8652 36654 8654 36706
rect 8706 36654 8708 36706
rect 8652 36642 8708 36654
rect 7980 36596 8036 36606
rect 7980 36502 8036 36540
rect 9100 36596 9156 36606
rect 9100 36502 9156 36540
rect 11228 36594 11284 36876
rect 11228 36542 11230 36594
rect 11282 36542 11284 36594
rect 11228 36530 11284 36542
rect 7812 35644 7924 35700
rect 8204 36482 8260 36494
rect 8204 36430 8206 36482
rect 8258 36430 8260 36482
rect 7756 35606 7812 35644
rect 7308 35534 7310 35586
rect 7362 35534 7364 35586
rect 7308 35522 7364 35534
rect 5180 35420 5796 35476
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 8204 34804 8260 36430
rect 12012 36484 12068 36494
rect 12460 36484 12516 36494
rect 12012 36482 12516 36484
rect 12012 36430 12014 36482
rect 12066 36430 12462 36482
rect 12514 36430 12516 36482
rect 12012 36428 12516 36430
rect 12012 36418 12068 36428
rect 12460 35700 12516 36428
rect 12460 35634 12516 35644
rect 13244 35700 13300 35710
rect 13244 35606 13300 35644
rect 13356 35028 13412 38108
rect 15036 38164 15092 40348
rect 15148 43538 15316 43540
rect 15148 43486 15262 43538
rect 15314 43486 15316 43538
rect 15148 43484 15316 43486
rect 15148 40290 15204 43484
rect 15260 43474 15316 43484
rect 15372 43484 15652 43540
rect 15372 42866 15428 43484
rect 15372 42814 15374 42866
rect 15426 42814 15428 42866
rect 15372 42802 15428 42814
rect 15484 43314 15540 43326
rect 15484 43262 15486 43314
rect 15538 43262 15540 43314
rect 15484 42868 15540 43262
rect 15596 43316 15652 43484
rect 15708 43538 15764 43652
rect 15708 43486 15710 43538
rect 15762 43486 15764 43538
rect 15708 43474 15764 43486
rect 18060 43540 18116 45388
rect 19964 45108 20020 45118
rect 20188 45108 20244 45388
rect 20636 45220 20692 45230
rect 20748 45220 20804 47182
rect 21980 46564 22036 47406
rect 23212 47458 23268 47628
rect 23212 47406 23214 47458
rect 23266 47406 23268 47458
rect 23212 47394 23268 47406
rect 23436 48244 23492 48254
rect 23436 47346 23492 48188
rect 24220 47458 24276 49532
rect 24780 49588 24836 49598
rect 24780 49494 24836 49532
rect 24892 49140 24948 49646
rect 25116 49700 25172 50430
rect 25900 50484 25956 50494
rect 25788 49924 25844 49934
rect 25788 49830 25844 49868
rect 25116 49634 25172 49644
rect 25676 49700 25732 49710
rect 25676 49606 25732 49644
rect 24892 49074 24948 49084
rect 25900 49028 25956 50428
rect 26236 50484 26292 51214
rect 27244 50706 27300 56030
rect 27804 55970 27860 56590
rect 49084 56642 49140 59200
rect 49084 56590 49086 56642
rect 49138 56590 49140 56642
rect 49084 56578 49140 56590
rect 49980 56642 50036 56654
rect 49980 56590 49982 56642
rect 50034 56590 50036 56642
rect 27804 55918 27806 55970
rect 27858 55918 27860 55970
rect 27804 55906 27860 55918
rect 49308 56082 49364 56094
rect 49308 56030 49310 56082
rect 49362 56030 49364 56082
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 49308 55468 49364 56030
rect 49980 55970 50036 56590
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 49980 55918 49982 55970
rect 50034 55918 50036 55970
rect 49980 55906 50036 55918
rect 48748 55412 49364 55468
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 41580 51492 41636 51502
rect 40796 51490 41636 51492
rect 40796 51438 41582 51490
rect 41634 51438 41636 51490
rect 40796 51436 41636 51438
rect 27244 50654 27246 50706
rect 27298 50654 27300 50706
rect 27244 50642 27300 50654
rect 33964 51378 34020 51390
rect 33964 51326 33966 51378
rect 34018 51326 34020 51378
rect 26236 50418 26292 50428
rect 27692 50484 27748 50494
rect 27692 50370 27748 50428
rect 27692 50318 27694 50370
rect 27746 50318 27748 50370
rect 27692 49810 27748 50318
rect 27692 49758 27694 49810
rect 27746 49758 27748 49810
rect 26460 49700 26516 49710
rect 26460 49606 26516 49644
rect 27132 49698 27188 49710
rect 27132 49646 27134 49698
rect 27186 49646 27188 49698
rect 25228 49026 25956 49028
rect 25228 48974 25902 49026
rect 25954 48974 25956 49026
rect 25228 48972 25956 48974
rect 25116 48916 25172 48926
rect 25116 48822 25172 48860
rect 25228 48692 25284 48972
rect 25900 48962 25956 48972
rect 26012 49586 26068 49598
rect 26012 49534 26014 49586
rect 26066 49534 26068 49586
rect 25116 48636 25284 48692
rect 24668 48468 24724 48478
rect 24668 48374 24724 48412
rect 24444 48356 24500 48366
rect 24444 48262 24500 48300
rect 24332 48244 24388 48254
rect 24332 48150 24388 48188
rect 24332 47572 24388 47582
rect 24332 47478 24388 47516
rect 24220 47406 24222 47458
rect 24274 47406 24276 47458
rect 24220 47394 24276 47406
rect 25116 47458 25172 48636
rect 25116 47406 25118 47458
rect 25170 47406 25172 47458
rect 25116 47394 25172 47406
rect 25564 48468 25620 48478
rect 23436 47294 23438 47346
rect 23490 47294 23492 47346
rect 23436 47124 23492 47294
rect 24108 47346 24164 47358
rect 24108 47294 24110 47346
rect 24162 47294 24164 47346
rect 23436 47068 23716 47124
rect 21980 46508 22260 46564
rect 21756 46116 21812 46126
rect 21756 46022 21812 46060
rect 20860 46004 20916 46014
rect 20860 45910 20916 45948
rect 21868 46004 21924 46014
rect 21868 45910 21924 45948
rect 22092 45890 22148 45902
rect 22092 45838 22094 45890
rect 22146 45838 22148 45890
rect 20636 45218 20804 45220
rect 20636 45166 20638 45218
rect 20690 45166 20804 45218
rect 20636 45164 20804 45166
rect 21644 45444 21700 45454
rect 20636 45154 20692 45164
rect 19964 45106 20244 45108
rect 19964 45054 19966 45106
rect 20018 45054 20244 45106
rect 19964 45052 20244 45054
rect 19964 45042 20020 45052
rect 19292 44098 19348 44110
rect 19292 44046 19294 44098
rect 19346 44046 19348 44098
rect 19292 43708 19348 44046
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19068 43652 19348 43708
rect 19068 43650 19124 43652
rect 19068 43598 19070 43650
rect 19122 43598 19124 43650
rect 19068 43586 19124 43598
rect 18060 43474 18116 43484
rect 18396 43540 18452 43550
rect 15932 43316 15988 43326
rect 15596 43314 15988 43316
rect 15596 43262 15934 43314
rect 15986 43262 15988 43314
rect 15596 43260 15988 43262
rect 15932 43250 15988 43260
rect 16044 43314 16100 43326
rect 16044 43262 16046 43314
rect 16098 43262 16100 43314
rect 16044 42980 16100 43262
rect 16044 42914 16100 42924
rect 15484 42802 15540 42812
rect 15148 40238 15150 40290
rect 15202 40238 15204 40290
rect 15148 40226 15204 40238
rect 15596 42756 15652 42766
rect 15036 38098 15092 38108
rect 14700 38052 14756 38062
rect 14700 37154 14756 37996
rect 15484 38052 15540 38062
rect 15484 37958 15540 37996
rect 15596 37826 15652 42700
rect 18284 42756 18340 42766
rect 18396 42756 18452 43484
rect 18844 43540 18900 43550
rect 18844 42866 18900 43484
rect 20188 43540 20244 45052
rect 20188 43474 20244 43484
rect 20860 44324 20916 44334
rect 18844 42814 18846 42866
rect 18898 42814 18900 42866
rect 18844 42802 18900 42814
rect 18284 42754 18452 42756
rect 18284 42702 18286 42754
rect 18338 42702 18452 42754
rect 18284 42700 18452 42702
rect 18284 42690 18340 42700
rect 17500 42642 17556 42654
rect 17500 42590 17502 42642
rect 17554 42590 17556 42642
rect 16492 42196 16548 42206
rect 16492 42102 16548 42140
rect 17500 42196 17556 42590
rect 20300 42532 20356 42542
rect 20188 42530 20356 42532
rect 20188 42478 20302 42530
rect 20354 42478 20356 42530
rect 20188 42476 20356 42478
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 17500 42130 17556 42140
rect 20188 42082 20244 42476
rect 20300 42466 20356 42476
rect 20860 42530 20916 44268
rect 21644 43650 21700 45388
rect 21756 44324 21812 44334
rect 21756 44230 21812 44268
rect 21644 43598 21646 43650
rect 21698 43598 21700 43650
rect 21644 43586 21700 43598
rect 21196 43428 21252 43438
rect 21196 43334 21252 43372
rect 22092 43428 22148 45838
rect 22204 45666 22260 46508
rect 22876 46562 22932 46574
rect 22876 46510 22878 46562
rect 22930 46510 22932 46562
rect 22876 46004 22932 46510
rect 22876 46002 23268 46004
rect 22876 45950 22878 46002
rect 22930 45950 23268 46002
rect 22876 45948 23268 45950
rect 22876 45938 22932 45948
rect 22316 45892 22372 45902
rect 22316 45890 22820 45892
rect 22316 45838 22318 45890
rect 22370 45838 22820 45890
rect 22316 45836 22820 45838
rect 22316 45826 22372 45836
rect 22204 45614 22206 45666
rect 22258 45614 22260 45666
rect 22204 45602 22260 45614
rect 22764 44994 22820 45836
rect 23212 45444 23268 45948
rect 23212 45330 23268 45388
rect 23212 45278 23214 45330
rect 23266 45278 23268 45330
rect 23212 45266 23268 45278
rect 22764 44942 22766 44994
rect 22818 44942 22820 44994
rect 22764 44930 22820 44942
rect 22540 44212 22596 44222
rect 22540 44118 22596 44156
rect 22092 43362 22148 43372
rect 23548 42868 23604 42878
rect 23548 42774 23604 42812
rect 20860 42478 20862 42530
rect 20914 42478 20916 42530
rect 20188 42030 20190 42082
rect 20242 42030 20244 42082
rect 20188 42018 20244 42030
rect 15820 41972 15876 41982
rect 15820 41878 15876 41916
rect 19404 41972 19460 41982
rect 17164 41188 17220 41198
rect 17164 39618 17220 41132
rect 17724 41188 17780 41198
rect 17724 41094 17780 41132
rect 19404 41188 19460 41916
rect 19404 41122 19460 41132
rect 20300 41972 20356 41982
rect 18508 41076 18564 41086
rect 18060 41074 18564 41076
rect 18060 41022 18510 41074
rect 18562 41022 18564 41074
rect 18060 41020 18564 41022
rect 18060 40626 18116 41020
rect 18508 41010 18564 41020
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 18060 40574 18062 40626
rect 18114 40574 18116 40626
rect 18060 40562 18116 40574
rect 19964 40516 20020 40526
rect 19068 40404 19124 40414
rect 19068 40310 19124 40348
rect 19964 39730 20020 40460
rect 19964 39678 19966 39730
rect 20018 39678 20020 39730
rect 19964 39666 20020 39678
rect 17164 39566 17166 39618
rect 17218 39566 17220 39618
rect 17164 39554 17220 39566
rect 17836 39506 17892 39518
rect 17836 39454 17838 39506
rect 17890 39454 17892 39506
rect 17836 39060 17892 39454
rect 20300 39396 20356 41916
rect 20860 41972 20916 42478
rect 20860 41906 20916 41916
rect 22316 41860 22372 41870
rect 22092 41858 22372 41860
rect 22092 41806 22318 41858
rect 22370 41806 22372 41858
rect 22092 41804 22372 41806
rect 22092 41410 22148 41804
rect 22316 41794 22372 41804
rect 22764 41858 22820 41870
rect 22764 41806 22766 41858
rect 22818 41806 22820 41858
rect 22092 41358 22094 41410
rect 22146 41358 22148 41410
rect 22092 41346 22148 41358
rect 20636 41300 20692 41310
rect 20636 41206 20692 41244
rect 21868 41300 21924 41310
rect 21868 41206 21924 41244
rect 21644 41186 21700 41198
rect 21644 41134 21646 41186
rect 21698 41134 21700 41186
rect 21644 40516 21700 41134
rect 21644 40450 21700 40460
rect 22316 41186 22372 41198
rect 22316 41134 22318 41186
rect 22370 41134 22372 41186
rect 21084 40404 21140 40414
rect 21084 40310 21140 40348
rect 22316 39844 22372 41134
rect 22428 41076 22484 41086
rect 22652 41076 22708 41086
rect 22428 41074 22708 41076
rect 22428 41022 22430 41074
rect 22482 41022 22654 41074
rect 22706 41022 22708 41074
rect 22428 41020 22708 41022
rect 22428 41010 22484 41020
rect 22652 41010 22708 41020
rect 22316 39788 22708 39844
rect 22316 39620 22372 39630
rect 22316 39526 22372 39564
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 17948 39060 18004 39070
rect 17836 39058 18004 39060
rect 17836 39006 17950 39058
rect 18002 39006 18004 39058
rect 17836 39004 18004 39006
rect 17948 38994 18004 39004
rect 20300 38834 20356 39340
rect 20860 39394 20916 39406
rect 20860 39342 20862 39394
rect 20914 39342 20916 39394
rect 20860 38948 20916 39342
rect 21532 39396 21588 39406
rect 21532 39302 21588 39340
rect 22652 39172 22708 39788
rect 22764 39396 22820 41806
rect 23660 41412 23716 47068
rect 24108 45332 24164 47294
rect 24668 46786 24724 46798
rect 24668 46734 24670 46786
rect 24722 46734 24724 46786
rect 24668 45892 24724 46734
rect 24780 46564 24836 46574
rect 25564 46564 25620 48412
rect 26012 48468 26068 49534
rect 26684 49588 26740 49598
rect 26012 48402 26068 48412
rect 26348 49026 26404 49038
rect 26348 48974 26350 49026
rect 26402 48974 26404 49026
rect 25676 48132 25732 48142
rect 25676 47572 25732 48076
rect 26348 48132 26404 48974
rect 26684 49026 26740 49532
rect 26684 48974 26686 49026
rect 26738 48974 26740 49026
rect 26684 48962 26740 48974
rect 26572 48916 26628 48926
rect 26572 48822 26628 48860
rect 27020 48916 27076 48926
rect 27132 48916 27188 49646
rect 27020 48914 27188 48916
rect 27020 48862 27022 48914
rect 27074 48862 27188 48914
rect 27020 48860 27188 48862
rect 27356 49700 27412 49710
rect 27020 48692 27076 48860
rect 27020 48626 27076 48636
rect 26348 48066 26404 48076
rect 27356 48242 27412 49644
rect 27356 48190 27358 48242
rect 27410 48190 27412 48242
rect 25788 48020 25844 48030
rect 25788 48018 26068 48020
rect 25788 47966 25790 48018
rect 25842 47966 26068 48018
rect 25788 47964 26068 47966
rect 25788 47954 25844 47964
rect 25732 47516 25956 47572
rect 25676 47440 25732 47516
rect 25788 47346 25844 47358
rect 25788 47294 25790 47346
rect 25842 47294 25844 47346
rect 25676 46788 25732 46798
rect 25788 46788 25844 47294
rect 25676 46786 25844 46788
rect 25676 46734 25678 46786
rect 25730 46734 25844 46786
rect 25676 46732 25844 46734
rect 25676 46722 25732 46732
rect 25788 46564 25844 46574
rect 25564 46562 25844 46564
rect 25564 46510 25790 46562
rect 25842 46510 25844 46562
rect 25564 46508 25844 46510
rect 24780 46470 24836 46508
rect 25788 46498 25844 46508
rect 24668 45826 24724 45836
rect 24892 46450 24948 46462
rect 24892 46398 24894 46450
rect 24946 46398 24948 46450
rect 24108 45266 24164 45276
rect 24668 44884 24724 44894
rect 24668 44434 24724 44828
rect 24892 44548 24948 46398
rect 25900 46114 25956 47516
rect 26012 46674 26068 47964
rect 26012 46622 26014 46674
rect 26066 46622 26068 46674
rect 26012 46610 26068 46622
rect 26908 46676 26964 46686
rect 26124 46564 26180 46574
rect 26124 46470 26180 46508
rect 26908 46562 26964 46620
rect 26908 46510 26910 46562
rect 26962 46510 26964 46562
rect 25900 46062 25902 46114
rect 25954 46062 25956 46114
rect 25900 46050 25956 46062
rect 25564 45890 25620 45902
rect 26124 45892 26180 45902
rect 25564 45838 25566 45890
rect 25618 45838 25620 45890
rect 25564 45220 25620 45838
rect 26012 45890 26180 45892
rect 26012 45838 26126 45890
rect 26178 45838 26180 45890
rect 26012 45836 26180 45838
rect 25564 45154 25620 45164
rect 25788 45778 25844 45790
rect 25788 45726 25790 45778
rect 25842 45726 25844 45778
rect 25788 45106 25844 45726
rect 26012 45332 26068 45836
rect 26124 45826 26180 45836
rect 26796 45892 26852 45902
rect 26796 45798 26852 45836
rect 26684 45332 26740 45342
rect 26908 45332 26964 46510
rect 26012 45276 26404 45332
rect 25788 45054 25790 45106
rect 25842 45054 25844 45106
rect 25788 44884 25844 45054
rect 25788 44818 25844 44828
rect 25900 45108 25956 45118
rect 24892 44482 24948 44492
rect 25452 44548 25508 44558
rect 25452 44454 25508 44492
rect 24668 44382 24670 44434
rect 24722 44382 24724 44434
rect 24668 44370 24724 44382
rect 25900 44322 25956 45052
rect 26012 45106 26068 45276
rect 26012 45054 26014 45106
rect 26066 45054 26068 45106
rect 26012 45042 26068 45054
rect 26236 45108 26292 45118
rect 26236 45014 26292 45052
rect 26124 44994 26180 45006
rect 26124 44942 26126 44994
rect 26178 44942 26180 44994
rect 25900 44270 25902 44322
rect 25954 44270 25956 44322
rect 25900 43538 25956 44270
rect 26012 44772 26068 44782
rect 26012 44322 26068 44716
rect 26124 44548 26180 44942
rect 26124 44482 26180 44492
rect 26012 44270 26014 44322
rect 26066 44270 26068 44322
rect 26012 44258 26068 44270
rect 26236 44324 26292 44334
rect 26348 44324 26404 45276
rect 26740 45276 27188 45332
rect 26684 45238 26740 45276
rect 26908 44660 26964 44670
rect 26908 44546 26964 44604
rect 26908 44494 26910 44546
rect 26962 44494 26964 44546
rect 26908 44482 26964 44494
rect 27132 44546 27188 45276
rect 27132 44494 27134 44546
rect 27186 44494 27188 44546
rect 27132 44482 27188 44494
rect 27244 44548 27300 44558
rect 27244 44454 27300 44492
rect 26236 44322 26404 44324
rect 26236 44270 26238 44322
rect 26290 44270 26404 44322
rect 26236 44268 26404 44270
rect 26236 43708 26292 44268
rect 26796 44212 26852 44222
rect 26796 44118 26852 44156
rect 25900 43486 25902 43538
rect 25954 43486 25956 43538
rect 25900 43474 25956 43486
rect 26124 43652 26292 43708
rect 26124 43538 26180 43652
rect 26124 43486 26126 43538
rect 26178 43486 26180 43538
rect 26012 43314 26068 43326
rect 26012 43262 26014 43314
rect 26066 43262 26068 43314
rect 25676 42642 25732 42654
rect 25676 42590 25678 42642
rect 25730 42590 25732 42642
rect 25676 41858 25732 42590
rect 25788 42196 25844 42206
rect 25788 42102 25844 42140
rect 26012 42082 26068 43262
rect 26124 42868 26180 43486
rect 26124 42802 26180 42812
rect 26012 42030 26014 42082
rect 26066 42030 26068 42082
rect 26012 42018 26068 42030
rect 26460 42754 26516 42766
rect 26460 42702 26462 42754
rect 26514 42702 26516 42754
rect 26460 41972 26516 42702
rect 26572 42196 26628 42206
rect 26572 42102 26628 42140
rect 26460 41906 26516 41916
rect 25676 41806 25678 41858
rect 25730 41806 25732 41858
rect 25676 41794 25732 41806
rect 23772 41412 23828 41422
rect 23660 41410 23828 41412
rect 23660 41358 23774 41410
rect 23826 41358 23828 41410
rect 23660 41356 23828 41358
rect 23772 41346 23828 41356
rect 22988 41186 23044 41198
rect 22988 41134 22990 41186
rect 23042 41134 23044 41186
rect 22876 41076 22932 41086
rect 22988 41076 23044 41134
rect 22876 41074 23044 41076
rect 22876 41022 22878 41074
rect 22930 41022 23044 41074
rect 22876 41020 23044 41022
rect 23212 41076 23268 41086
rect 22876 41010 22932 41020
rect 23212 40982 23268 41020
rect 23324 41074 23380 41086
rect 23324 41022 23326 41074
rect 23378 41022 23380 41074
rect 22988 40516 23044 40526
rect 22988 39730 23044 40460
rect 22988 39678 22990 39730
rect 23042 39678 23044 39730
rect 22988 39666 23044 39678
rect 22764 39330 22820 39340
rect 22652 39116 23156 39172
rect 20972 38948 21028 38958
rect 20860 38946 21028 38948
rect 20860 38894 20974 38946
rect 21026 38894 21028 38946
rect 20860 38892 21028 38894
rect 20972 38882 21028 38892
rect 20300 38782 20302 38834
rect 20354 38782 20356 38834
rect 20300 38770 20356 38782
rect 15708 38722 15764 38734
rect 15708 38670 15710 38722
rect 15762 38670 15764 38722
rect 15708 38274 15764 38670
rect 23100 38722 23156 39116
rect 23100 38670 23102 38722
rect 23154 38670 23156 38722
rect 23100 38658 23156 38670
rect 15708 38222 15710 38274
rect 15762 38222 15764 38274
rect 15708 38210 15764 38222
rect 15932 38052 15988 38062
rect 15932 38050 16100 38052
rect 15932 37998 15934 38050
rect 15986 37998 16100 38050
rect 15932 37996 16100 37998
rect 15932 37986 15988 37996
rect 15596 37774 15598 37826
rect 15650 37774 15652 37826
rect 15596 37762 15652 37774
rect 15932 37380 15988 37390
rect 14700 37102 14702 37154
rect 14754 37102 14756 37154
rect 14700 37090 14756 37102
rect 15260 37378 15988 37380
rect 15260 37326 15934 37378
rect 15986 37326 15988 37378
rect 15260 37324 15988 37326
rect 15260 36594 15316 37324
rect 15932 37314 15988 37324
rect 15260 36542 15262 36594
rect 15314 36542 15316 36594
rect 15260 36530 15316 36542
rect 14476 36482 14532 36494
rect 14476 36430 14478 36482
rect 14530 36430 14532 36482
rect 13916 36258 13972 36270
rect 13916 36206 13918 36258
rect 13970 36206 13972 36258
rect 13916 35812 13972 36206
rect 14028 35812 14084 35822
rect 13916 35810 14084 35812
rect 13916 35758 14030 35810
rect 14082 35758 14084 35810
rect 13916 35756 14084 35758
rect 14028 35746 14084 35756
rect 14476 35700 14532 36430
rect 14476 35634 14532 35644
rect 16044 35588 16100 37996
rect 16156 38050 16212 38062
rect 16156 37998 16158 38050
rect 16210 37998 16212 38050
rect 16156 36596 16212 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 17724 37154 17780 37166
rect 17724 37102 17726 37154
rect 17778 37102 17780 37154
rect 16156 36530 16212 36540
rect 17388 36596 17444 36606
rect 17388 36502 17444 36540
rect 17724 36484 17780 37102
rect 20860 36594 20916 36606
rect 20860 36542 20862 36594
rect 20914 36542 20916 36594
rect 17948 36484 18004 36494
rect 17724 36482 18004 36484
rect 17724 36430 17950 36482
rect 18002 36430 18004 36482
rect 17724 36428 18004 36430
rect 16604 35700 16660 35710
rect 17612 35700 17668 35710
rect 16660 35644 16884 35700
rect 16604 35606 16660 35644
rect 16156 35588 16212 35598
rect 16044 35586 16212 35588
rect 16044 35534 16158 35586
rect 16210 35534 16212 35586
rect 16044 35532 16212 35534
rect 16156 35522 16212 35532
rect 13692 35028 13748 35038
rect 13356 35026 13748 35028
rect 13356 34974 13694 35026
rect 13746 34974 13748 35026
rect 13356 34972 13748 34974
rect 13692 34916 13748 34972
rect 16828 35028 16884 35644
rect 17612 35606 17668 35644
rect 17948 35700 18004 36428
rect 18732 36372 18788 36382
rect 18732 36370 19684 36372
rect 18732 36318 18734 36370
rect 18786 36318 19684 36370
rect 18732 36316 19684 36318
rect 18732 36306 18788 36316
rect 19628 35924 19684 36316
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19740 35924 19796 35934
rect 19628 35922 19796 35924
rect 19628 35870 19742 35922
rect 19794 35870 19796 35922
rect 19628 35868 19796 35870
rect 19740 35858 19796 35868
rect 18844 35812 18900 35822
rect 18620 35810 18900 35812
rect 18620 35758 18846 35810
rect 18898 35758 18900 35810
rect 18620 35756 18900 35758
rect 17948 35634 18004 35644
rect 18284 35700 18340 35710
rect 16828 35026 17220 35028
rect 16828 34974 16830 35026
rect 16882 34974 17220 35026
rect 16828 34972 17220 34974
rect 16828 34962 16884 34972
rect 8204 34738 8260 34748
rect 8988 34804 9044 34814
rect 6188 34130 6244 34142
rect 6188 34078 6190 34130
rect 6242 34078 6244 34130
rect 6188 34020 6244 34078
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 5964 31108 6020 31118
rect 5964 30994 6020 31052
rect 6188 31108 6244 33964
rect 6860 34020 6916 34030
rect 6860 34018 7140 34020
rect 6860 33966 6862 34018
rect 6914 33966 7140 34018
rect 6860 33964 7140 33966
rect 6860 33954 6916 33964
rect 7084 33234 7140 33964
rect 8988 34018 9044 34748
rect 13692 34242 13748 34860
rect 14252 34916 14308 34926
rect 14252 34822 14308 34860
rect 15036 34916 15092 34926
rect 13692 34190 13694 34242
rect 13746 34190 13748 34242
rect 13692 34178 13748 34190
rect 8988 33966 8990 34018
rect 9042 33966 9044 34018
rect 8988 33954 9044 33966
rect 9772 34020 9828 34030
rect 9772 33926 9828 33964
rect 12236 34020 12292 34030
rect 7084 33182 7086 33234
rect 7138 33182 7140 33234
rect 7084 33170 7140 33182
rect 11228 33122 11284 33134
rect 11228 33070 11230 33122
rect 11282 33070 11284 33122
rect 11228 31948 11284 33070
rect 10780 31892 11284 31948
rect 12236 32786 12292 33964
rect 14364 33458 14420 33470
rect 14364 33406 14366 33458
rect 14418 33406 14420 33458
rect 13692 33122 13748 33134
rect 13692 33070 13694 33122
rect 13746 33070 13748 33122
rect 12236 32734 12238 32786
rect 12290 32734 12292 32786
rect 10780 31890 10836 31892
rect 10780 31838 10782 31890
rect 10834 31838 10836 31890
rect 10780 31826 10836 31838
rect 10108 31778 10164 31790
rect 10108 31726 10110 31778
rect 10162 31726 10164 31778
rect 6188 31042 6244 31052
rect 6412 31108 6468 31118
rect 6412 31014 6468 31052
rect 10108 31108 10164 31726
rect 5964 30942 5966 30994
rect 6018 30942 6020 30994
rect 5964 30930 6020 30942
rect 5068 30884 5124 30894
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5068 29540 5124 30828
rect 5180 30882 5236 30894
rect 5180 30830 5182 30882
rect 5234 30830 5236 30882
rect 5180 30436 5236 30830
rect 5180 30380 6020 30436
rect 5852 30212 5908 30222
rect 5516 30210 5908 30212
rect 5516 30158 5854 30210
rect 5906 30158 5908 30210
rect 5516 30156 5908 30158
rect 5180 29540 5236 29550
rect 5068 29538 5236 29540
rect 5068 29486 5182 29538
rect 5234 29486 5236 29538
rect 5068 29484 5236 29486
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4172 28690 4228 28700
rect 5180 28644 5236 29484
rect 5180 28578 5236 28588
rect 5404 29538 5460 29550
rect 5404 29486 5406 29538
rect 5458 29486 5460 29538
rect 5404 28532 5460 29486
rect 5516 29314 5572 30156
rect 5852 30146 5908 30156
rect 5964 29986 6020 30380
rect 6076 30212 6132 30222
rect 6300 30212 6356 30222
rect 10108 30212 10164 31052
rect 6076 30210 6244 30212
rect 6076 30158 6078 30210
rect 6130 30158 6244 30210
rect 6076 30156 6244 30158
rect 6076 30146 6132 30156
rect 5964 29934 5966 29986
rect 6018 29934 6020 29986
rect 5964 29922 6020 29934
rect 6076 29316 6132 29326
rect 5516 29262 5518 29314
rect 5570 29262 5572 29314
rect 5516 29250 5572 29262
rect 5964 29314 6132 29316
rect 5964 29262 6078 29314
rect 6130 29262 6132 29314
rect 5964 29260 6132 29262
rect 5404 28466 5460 28476
rect 5964 28642 6020 29260
rect 6076 29250 6132 29260
rect 6188 28980 6244 30156
rect 6300 30210 6692 30212
rect 6300 30158 6302 30210
rect 6354 30158 6692 30210
rect 6300 30156 6692 30158
rect 6300 30146 6356 30156
rect 5964 28590 5966 28642
rect 6018 28590 6020 28642
rect 5964 28532 6020 28590
rect 5964 28466 6020 28476
rect 6076 28924 6580 28980
rect 6076 27970 6132 28924
rect 6524 28866 6580 28924
rect 6524 28814 6526 28866
rect 6578 28814 6580 28866
rect 6188 28644 6244 28654
rect 6188 28550 6244 28588
rect 6076 27918 6078 27970
rect 6130 27918 6132 27970
rect 6076 27906 6132 27918
rect 6300 27970 6356 27982
rect 6300 27918 6302 27970
rect 6354 27918 6356 27970
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 6300 27186 6356 27918
rect 6300 27134 6302 27186
rect 6354 27134 6356 27186
rect 3388 26290 3444 26302
rect 3388 26238 3390 26290
rect 3442 26238 3444 26290
rect 2716 23492 2772 23502
rect 2716 23154 2772 23436
rect 3388 23492 3444 26238
rect 4172 26180 4228 26190
rect 4172 26086 4228 26124
rect 6188 26180 6244 26190
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 6188 25730 6244 26124
rect 6300 26178 6356 27134
rect 6412 27634 6468 27646
rect 6412 27582 6414 27634
rect 6466 27582 6468 27634
rect 6412 27076 6468 27582
rect 6524 27298 6580 28814
rect 6636 28868 6692 30156
rect 9660 30156 10164 30212
rect 9660 29650 9716 30156
rect 9660 29598 9662 29650
rect 9714 29598 9716 29650
rect 8988 29428 9044 29438
rect 8988 29334 9044 29372
rect 9660 29428 9716 29598
rect 9660 29362 9716 29372
rect 8204 29316 8260 29326
rect 6636 28802 6692 28812
rect 7420 29314 8260 29316
rect 7420 29262 8206 29314
rect 8258 29262 8260 29314
rect 7420 29260 8260 29262
rect 7420 28754 7476 29260
rect 8204 29250 8260 29260
rect 7532 28868 7588 28878
rect 7532 28774 7588 28812
rect 8204 28868 8260 28878
rect 7420 28702 7422 28754
rect 7474 28702 7476 28754
rect 7420 28690 7476 28702
rect 7308 28532 7364 28542
rect 7308 28438 7364 28476
rect 6524 27246 6526 27298
rect 6578 27246 6580 27298
rect 6524 27234 6580 27246
rect 6412 27020 6692 27076
rect 6300 26126 6302 26178
rect 6354 26126 6356 26178
rect 6300 26114 6356 26126
rect 6524 26852 6580 26862
rect 6188 25678 6190 25730
rect 6242 25678 6244 25730
rect 6188 25666 6244 25678
rect 6300 25732 6356 25742
rect 6300 25638 6356 25676
rect 6524 25730 6580 26796
rect 6524 25678 6526 25730
rect 6578 25678 6580 25730
rect 6524 25666 6580 25678
rect 6636 25730 6692 27020
rect 6860 26852 6916 26862
rect 6860 26758 6916 26796
rect 7532 26852 7588 26862
rect 7308 26404 7364 26414
rect 7308 26290 7364 26348
rect 7308 26238 7310 26290
rect 7362 26238 7364 26290
rect 6636 25678 6638 25730
rect 6690 25678 6692 25730
rect 6636 25666 6692 25678
rect 6860 26178 6916 26190
rect 6860 26126 6862 26178
rect 6914 26126 6916 26178
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4620 23716 4676 23726
rect 3388 23426 3444 23436
rect 3500 23714 4676 23716
rect 3500 23662 4622 23714
rect 4674 23662 4676 23714
rect 3500 23660 4676 23662
rect 3388 23268 3444 23278
rect 3500 23268 3556 23660
rect 4620 23650 4676 23660
rect 5740 23714 5796 23726
rect 5740 23662 5742 23714
rect 5794 23662 5796 23714
rect 3388 23266 3556 23268
rect 3388 23214 3390 23266
rect 3442 23214 3556 23266
rect 3388 23212 3556 23214
rect 3948 23492 4004 23502
rect 3388 23202 3444 23212
rect 2716 23102 2718 23154
rect 2770 23102 2772 23154
rect 1820 22482 1876 22494
rect 1820 22430 1822 22482
rect 1874 22430 1876 22482
rect 1820 21586 1876 22430
rect 1820 21534 1822 21586
rect 1874 21534 1876 21586
rect 1820 21522 1876 21534
rect 2268 21924 2324 21934
rect 2268 20188 2324 21868
rect 2716 21924 2772 23102
rect 3948 22482 4004 23436
rect 5740 23156 5796 23662
rect 6076 23268 6132 23278
rect 6076 23156 6132 23212
rect 6860 23268 6916 26126
rect 6972 25732 7028 25742
rect 6972 24834 7028 25676
rect 6972 24782 6974 24834
rect 7026 24782 7028 24834
rect 6972 24770 7028 24782
rect 7308 24722 7364 26238
rect 7532 26290 7588 26796
rect 8204 26850 8260 28812
rect 9996 28642 10052 30156
rect 12236 29652 12292 32734
rect 12908 32788 12964 32798
rect 12908 32562 12964 32732
rect 13580 32676 13636 32686
rect 13692 32676 13748 33070
rect 13580 32674 13748 32676
rect 13580 32622 13582 32674
rect 13634 32622 13748 32674
rect 13580 32620 13748 32622
rect 13804 32788 13860 32798
rect 13580 32610 13636 32620
rect 12908 32510 12910 32562
rect 12962 32510 12964 32562
rect 12908 32498 12964 32510
rect 12908 31890 12964 31902
rect 12908 31838 12910 31890
rect 12962 31838 12964 31890
rect 12908 31220 12964 31838
rect 13804 31778 13860 32732
rect 14364 31892 14420 33406
rect 14364 31826 14420 31836
rect 13804 31726 13806 31778
rect 13858 31726 13860 31778
rect 13804 31714 13860 31726
rect 14476 31668 14532 31678
rect 12908 31154 12964 31164
rect 13916 31666 14532 31668
rect 13916 31614 14478 31666
rect 14530 31614 14532 31666
rect 13916 31612 14532 31614
rect 13916 30098 13972 31612
rect 14476 31602 14532 31612
rect 15036 30996 15092 34860
rect 16492 34244 16548 34254
rect 15484 34132 15540 34142
rect 15036 30902 15092 30940
rect 15372 30996 15428 31006
rect 15372 30210 15428 30940
rect 15372 30158 15374 30210
rect 15426 30158 15428 30210
rect 15372 30146 15428 30158
rect 13916 30046 13918 30098
rect 13970 30046 13972 30098
rect 13916 30034 13972 30046
rect 12236 29586 12292 29596
rect 13132 29652 13188 29662
rect 13132 29558 13188 29596
rect 11564 29540 11620 29550
rect 10780 29538 11620 29540
rect 10780 29486 11566 29538
rect 11618 29486 11620 29538
rect 10780 29484 11620 29486
rect 10780 28754 10836 29484
rect 11564 29474 11620 29484
rect 10780 28702 10782 28754
rect 10834 28702 10836 28754
rect 10780 28690 10836 28702
rect 12908 28754 12964 28766
rect 12908 28702 12910 28754
rect 12962 28702 12964 28754
rect 9996 28590 9998 28642
rect 10050 28590 10052 28642
rect 9996 28578 10052 28590
rect 9436 28420 9492 28430
rect 8988 27188 9044 27198
rect 9436 27188 9492 28364
rect 12908 27412 12964 28702
rect 15484 28644 15540 34076
rect 16492 33458 16548 34188
rect 16716 34132 16772 34142
rect 16716 34038 16772 34076
rect 16492 33406 16494 33458
rect 16546 33406 16548 33458
rect 16492 33394 16548 33406
rect 17164 33346 17220 34972
rect 18284 34354 18340 35644
rect 18284 34302 18286 34354
rect 18338 34302 18340 34354
rect 18284 34290 18340 34302
rect 17724 34244 17780 34254
rect 17724 34150 17780 34188
rect 18620 33458 18676 35756
rect 18844 35746 18900 35756
rect 20860 35140 20916 36542
rect 21980 36258 22036 36270
rect 21980 36206 21982 36258
rect 22034 36206 22036 36258
rect 21868 35812 21924 35822
rect 21980 35812 22036 36206
rect 21868 35810 22036 35812
rect 21868 35758 21870 35810
rect 21922 35758 22036 35810
rect 21868 35756 22036 35758
rect 21868 35746 21924 35756
rect 21196 35700 21252 35710
rect 21196 35606 21252 35644
rect 22988 35588 23044 35598
rect 20860 35074 20916 35084
rect 22428 35140 22484 35150
rect 22428 35046 22484 35084
rect 22988 35138 23044 35532
rect 22988 35086 22990 35138
rect 23042 35086 23044 35138
rect 22988 35074 23044 35086
rect 23100 35140 23156 35150
rect 23324 35140 23380 41022
rect 26908 41076 26964 41086
rect 24332 40962 24388 40974
rect 24332 40910 24334 40962
rect 24386 40910 24388 40962
rect 24332 40516 24388 40910
rect 24332 40450 24388 40460
rect 25676 40404 25732 40414
rect 25564 40402 25732 40404
rect 25564 40350 25678 40402
rect 25730 40350 25732 40402
rect 25564 40348 25732 40350
rect 23548 40290 23604 40302
rect 23548 40238 23550 40290
rect 23602 40238 23604 40290
rect 23548 39396 23604 40238
rect 25116 39730 25172 39742
rect 25116 39678 25118 39730
rect 25170 39678 25172 39730
rect 23548 38722 23604 39340
rect 23548 38670 23550 38722
rect 23602 38670 23604 38722
rect 23548 35700 23604 38670
rect 24556 39620 24612 39630
rect 24556 38050 24612 39564
rect 25116 38836 25172 39678
rect 25564 39620 25620 40348
rect 25676 40338 25732 40348
rect 26684 40404 26740 40414
rect 25676 39732 25732 39742
rect 25676 39638 25732 39676
rect 25564 39554 25620 39564
rect 25676 38948 25732 38958
rect 25116 38770 25172 38780
rect 25340 38946 25732 38948
rect 25340 38894 25678 38946
rect 25730 38894 25732 38946
rect 25340 38892 25732 38894
rect 25340 38162 25396 38892
rect 25676 38882 25732 38892
rect 25340 38110 25342 38162
rect 25394 38110 25396 38162
rect 25340 38098 25396 38110
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 24220 37492 24276 37502
rect 24220 37398 24276 37436
rect 24556 36484 24612 37998
rect 26684 37492 26740 40348
rect 26908 39058 26964 41020
rect 27020 40964 27076 40974
rect 27020 40962 27188 40964
rect 27020 40910 27022 40962
rect 27074 40910 27188 40962
rect 27020 40908 27188 40910
rect 27020 40898 27076 40908
rect 27132 40180 27188 40908
rect 27244 40404 27300 40414
rect 27356 40404 27412 48190
rect 27468 46676 27524 46686
rect 27468 46582 27524 46620
rect 27692 46676 27748 49758
rect 33964 50484 34020 51326
rect 34748 51266 34804 51278
rect 34748 51214 34750 51266
rect 34802 51214 34804 51266
rect 34748 50484 34804 51214
rect 36876 51268 36932 51278
rect 36876 51266 37380 51268
rect 36876 51214 36878 51266
rect 36930 51214 37380 51266
rect 36876 51212 37380 51214
rect 36876 51202 36932 51212
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 34860 50484 34916 50494
rect 34748 50482 34916 50484
rect 34748 50430 34862 50482
rect 34914 50430 34916 50482
rect 34748 50428 34916 50430
rect 28364 49698 28420 49710
rect 28364 49646 28366 49698
rect 28418 49646 28420 49698
rect 28364 49250 28420 49646
rect 28364 49198 28366 49250
rect 28418 49198 28420 49250
rect 28364 49186 28420 49198
rect 30492 49698 30548 49710
rect 30492 49646 30494 49698
rect 30546 49646 30548 49698
rect 30268 49026 30324 49038
rect 30268 48974 30270 49026
rect 30322 48974 30324 49026
rect 28700 48916 28756 48926
rect 28700 48822 28756 48860
rect 30044 48916 30100 48926
rect 30044 48822 30100 48860
rect 27692 46610 27748 46620
rect 27804 48802 27860 48814
rect 27804 48750 27806 48802
rect 27858 48750 27860 48802
rect 27804 48692 27860 48750
rect 27804 47348 27860 48636
rect 28476 48802 28532 48814
rect 28476 48750 28478 48802
rect 28530 48750 28532 48802
rect 27804 46786 27860 47292
rect 27804 46734 27806 46786
rect 27858 46734 27860 46786
rect 27804 42196 27860 46734
rect 27916 47570 27972 47582
rect 27916 47518 27918 47570
rect 27970 47518 27972 47570
rect 27916 45892 27972 47518
rect 28476 47348 28532 48750
rect 28812 47572 28868 47582
rect 28812 47570 29204 47572
rect 28812 47518 28814 47570
rect 28866 47518 29204 47570
rect 28812 47516 29204 47518
rect 28812 47506 28868 47516
rect 28476 47254 28532 47292
rect 28700 47460 28756 47470
rect 28700 47346 28756 47404
rect 28700 47294 28702 47346
rect 28754 47294 28756 47346
rect 28700 47282 28756 47294
rect 29148 46786 29204 47516
rect 30268 47460 30324 48974
rect 30492 49028 30548 49646
rect 30940 49700 30996 49710
rect 30940 49698 31108 49700
rect 30940 49646 30942 49698
rect 30994 49646 31108 49698
rect 30940 49644 31108 49646
rect 30940 49634 30996 49644
rect 30940 49028 30996 49038
rect 30492 49026 30996 49028
rect 30492 48974 30942 49026
rect 30994 48974 30996 49026
rect 30492 48972 30996 48974
rect 30268 47394 30324 47404
rect 30716 47460 30772 47470
rect 30716 47366 30772 47404
rect 29484 47348 29540 47358
rect 29484 47254 29540 47292
rect 30828 47348 30884 47358
rect 30940 47348 30996 48972
rect 31052 48132 31108 49644
rect 33852 48804 33908 48814
rect 33852 48710 33908 48748
rect 32508 48354 32564 48366
rect 32508 48302 32510 48354
rect 32562 48302 32564 48354
rect 31724 48132 31780 48142
rect 31052 48130 31780 48132
rect 31052 48078 31726 48130
rect 31778 48078 31780 48130
rect 31052 48076 31780 48078
rect 31052 47460 31108 47470
rect 31612 47460 31668 47470
rect 31052 47458 31668 47460
rect 31052 47406 31054 47458
rect 31106 47406 31614 47458
rect 31666 47406 31668 47458
rect 31052 47404 31668 47406
rect 31052 47394 31108 47404
rect 30828 47346 30940 47348
rect 30828 47294 30830 47346
rect 30882 47294 30940 47346
rect 30828 47292 30940 47294
rect 30828 47282 30884 47292
rect 29148 46734 29150 46786
rect 29202 46734 29204 46786
rect 29148 46722 29204 46734
rect 29820 47236 29876 47246
rect 27916 45826 27972 45836
rect 28476 46676 28532 46686
rect 28140 45666 28196 45678
rect 28140 45614 28142 45666
rect 28194 45614 28196 45666
rect 27916 45444 27972 45454
rect 27916 43538 27972 45388
rect 28140 45444 28196 45614
rect 28140 45378 28196 45388
rect 28476 45444 28532 46620
rect 29820 46114 29876 47180
rect 30268 47234 30324 47246
rect 30268 47182 30270 47234
rect 30322 47182 30324 47234
rect 29820 46062 29822 46114
rect 29874 46062 29876 46114
rect 29820 46050 29876 46062
rect 30156 46116 30212 46126
rect 30268 46116 30324 47182
rect 30156 46114 30772 46116
rect 30156 46062 30158 46114
rect 30210 46062 30772 46114
rect 30156 46060 30772 46062
rect 30156 46050 30212 46060
rect 29932 45890 29988 45902
rect 29932 45838 29934 45890
rect 29986 45838 29988 45890
rect 28476 45378 28532 45388
rect 28812 45666 28868 45678
rect 28812 45614 28814 45666
rect 28866 45614 28868 45666
rect 28812 45332 28868 45614
rect 29820 45668 29876 45678
rect 29820 45574 29876 45612
rect 28364 45218 28420 45230
rect 28364 45166 28366 45218
rect 28418 45166 28420 45218
rect 28140 45108 28196 45118
rect 28140 45014 28196 45052
rect 28364 44996 28420 45166
rect 28364 44930 28420 44940
rect 28812 44436 28868 45276
rect 29708 44996 29764 45006
rect 29708 44546 29764 44940
rect 29708 44494 29710 44546
rect 29762 44494 29764 44546
rect 29708 44482 29764 44494
rect 28924 44436 28980 44446
rect 28812 44380 28924 44436
rect 28924 44304 28980 44380
rect 29932 44436 29988 45838
rect 30604 45556 30660 45566
rect 30268 45108 30324 45118
rect 30268 45014 30324 45052
rect 30604 45106 30660 45500
rect 30604 45054 30606 45106
rect 30658 45054 30660 45106
rect 30604 45042 30660 45054
rect 30716 44546 30772 46060
rect 30828 46004 30884 46014
rect 30828 45910 30884 45948
rect 30940 45218 30996 47292
rect 31164 46228 31220 47404
rect 31612 47394 31668 47404
rect 31276 46564 31332 46574
rect 31332 46508 31444 46564
rect 31276 46470 31332 46508
rect 31164 46172 31332 46228
rect 31276 46004 31332 46172
rect 30940 45166 30942 45218
rect 30994 45166 30996 45218
rect 30940 45154 30996 45166
rect 31164 45444 31220 45454
rect 30716 44494 30718 44546
rect 30770 44494 30772 44546
rect 30716 44482 30772 44494
rect 31052 45106 31108 45118
rect 31052 45054 31054 45106
rect 31106 45054 31108 45106
rect 29932 44342 29988 44380
rect 30156 44324 30212 44334
rect 30156 44230 30212 44268
rect 30828 44324 30884 44334
rect 31052 44324 31108 45054
rect 30828 44230 30884 44268
rect 30940 44322 31108 44324
rect 30940 44270 31054 44322
rect 31106 44270 31108 44322
rect 30940 44268 31108 44270
rect 29596 44212 29652 44222
rect 29036 44210 29652 44212
rect 29036 44158 29598 44210
rect 29650 44158 29652 44210
rect 29036 44156 29652 44158
rect 29036 43764 29092 44156
rect 29596 44146 29652 44156
rect 30940 43988 30996 44268
rect 31052 44258 31108 44268
rect 28588 43708 29092 43764
rect 30716 43932 30996 43988
rect 28588 43650 28644 43708
rect 28588 43598 28590 43650
rect 28642 43598 28644 43650
rect 28588 43586 28644 43598
rect 27916 43486 27918 43538
rect 27970 43486 27972 43538
rect 27916 43474 27972 43486
rect 30716 43426 30772 43932
rect 31164 43762 31220 45388
rect 31276 45106 31332 45948
rect 31388 45556 31444 46508
rect 31388 45490 31444 45500
rect 31724 46562 31780 48076
rect 32172 47460 32228 47470
rect 32172 47366 32228 47404
rect 32508 47460 32564 48302
rect 32508 47394 32564 47404
rect 32732 48242 32788 48254
rect 32732 48190 32734 48242
rect 32786 48190 32788 48242
rect 31836 47348 31892 47358
rect 31836 47254 31892 47292
rect 31948 47236 32004 47246
rect 31948 47142 32004 47180
rect 31724 46510 31726 46562
rect 31778 46510 31780 46562
rect 31724 45444 31780 46510
rect 32732 46564 32788 48190
rect 33740 48244 33796 48254
rect 33964 48244 34020 50428
rect 34860 50418 34916 50428
rect 36316 50484 36372 50494
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 36316 49140 36372 50428
rect 36876 49812 36932 49822
rect 36876 49718 36932 49756
rect 36764 49140 36820 49150
rect 36316 49138 37044 49140
rect 36316 49086 36318 49138
rect 36370 49086 36766 49138
rect 36818 49086 37044 49138
rect 36316 49084 37044 49086
rect 36316 49074 36372 49084
rect 36764 49074 36820 49084
rect 34412 48804 34468 48814
rect 35196 48804 35252 48814
rect 34412 48354 34468 48748
rect 34412 48302 34414 48354
rect 34466 48302 34468 48354
rect 34412 48290 34468 48302
rect 34636 48802 35252 48804
rect 34636 48750 35198 48802
rect 35250 48750 35252 48802
rect 34636 48748 35252 48750
rect 33740 48242 34020 48244
rect 33740 48190 33742 48242
rect 33794 48190 34020 48242
rect 33740 48188 34020 48190
rect 33740 48178 33796 48188
rect 33852 47458 33908 48188
rect 34636 47570 34692 48748
rect 35196 48738 35252 48748
rect 36988 48468 37044 49084
rect 36988 48466 37156 48468
rect 36988 48414 36990 48466
rect 37042 48414 37156 48466
rect 36988 48412 37156 48414
rect 36988 48402 37044 48412
rect 36540 48130 36596 48142
rect 36540 48078 36542 48130
rect 36594 48078 36596 48130
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 36540 47684 36596 48078
rect 36540 47618 36596 47628
rect 34636 47518 34638 47570
rect 34690 47518 34692 47570
rect 34636 47506 34692 47518
rect 36764 47572 36820 47582
rect 36764 47478 36820 47516
rect 33852 47406 33854 47458
rect 33906 47406 33908 47458
rect 33852 47394 33908 47406
rect 37100 46898 37156 48412
rect 37324 47460 37380 51212
rect 37436 51266 37492 51278
rect 37436 51214 37438 51266
rect 37490 51214 37492 51266
rect 37436 50484 37492 51214
rect 40796 50706 40852 51436
rect 41580 51426 41636 51436
rect 45948 51378 46004 51390
rect 45948 51326 45950 51378
rect 46002 51326 46004 51378
rect 40796 50654 40798 50706
rect 40850 50654 40852 50706
rect 40796 50642 40852 50654
rect 42924 50706 42980 50718
rect 42924 50654 42926 50706
rect 42978 50654 42980 50706
rect 40012 50594 40068 50606
rect 40012 50542 40014 50594
rect 40066 50542 40068 50594
rect 39452 50484 39508 50494
rect 37492 50428 37604 50484
rect 37436 50418 37492 50428
rect 37548 49700 37604 50428
rect 39452 50390 39508 50428
rect 40012 50484 40068 50542
rect 40012 50418 40068 50428
rect 40348 50484 40404 50494
rect 37660 50372 37716 50382
rect 37660 50278 37716 50316
rect 39676 50372 39732 50382
rect 37884 49700 37940 49710
rect 37548 49698 37940 49700
rect 37548 49646 37886 49698
rect 37938 49646 37940 49698
rect 37548 49644 37940 49646
rect 37548 49140 37604 49150
rect 37548 49138 37828 49140
rect 37548 49086 37550 49138
rect 37602 49086 37828 49138
rect 37548 49084 37828 49086
rect 37548 49074 37604 49084
rect 37772 48020 37828 49084
rect 37884 48242 37940 49644
rect 39676 49138 39732 50316
rect 39676 49086 39678 49138
rect 39730 49086 39732 49138
rect 39676 49074 39732 49086
rect 40348 49028 40404 50428
rect 42700 50034 42756 50046
rect 42700 49982 42702 50034
rect 42754 49982 42756 50034
rect 41692 49922 41748 49934
rect 41692 49870 41694 49922
rect 41746 49870 41748 49922
rect 41692 49140 41748 49870
rect 42252 49812 42308 49822
rect 42140 49756 42252 49812
rect 41804 49140 41860 49150
rect 41692 49138 41860 49140
rect 41692 49086 41806 49138
rect 41858 49086 41860 49138
rect 41692 49084 41860 49086
rect 41804 49074 41860 49084
rect 41020 49028 41076 49038
rect 40348 49026 41524 49028
rect 40348 48974 40350 49026
rect 40402 48974 41022 49026
rect 41074 48974 41524 49026
rect 40348 48972 41524 48974
rect 40348 48962 40404 48972
rect 41020 48962 41076 48972
rect 41468 48466 41524 48972
rect 41468 48414 41470 48466
rect 41522 48414 41524 48466
rect 41468 48402 41524 48414
rect 37884 48190 37886 48242
rect 37938 48190 37940 48242
rect 37884 48178 37940 48190
rect 38668 48132 38724 48142
rect 40796 48132 40852 48142
rect 38668 48130 39172 48132
rect 38668 48078 38670 48130
rect 38722 48078 39172 48130
rect 38668 48076 39172 48078
rect 38668 48066 38724 48076
rect 37772 47964 38276 48020
rect 37772 47684 37828 47694
rect 37772 47590 37828 47628
rect 38220 47682 38276 47964
rect 38220 47630 38222 47682
rect 38274 47630 38276 47682
rect 38220 47618 38276 47630
rect 37996 47572 38052 47582
rect 37996 47478 38052 47516
rect 37548 47460 37604 47470
rect 37324 47458 37604 47460
rect 37324 47406 37550 47458
rect 37602 47406 37604 47458
rect 37324 47404 37604 47406
rect 37548 47394 37604 47404
rect 38332 47346 38388 47358
rect 38332 47294 38334 47346
rect 38386 47294 38388 47346
rect 38332 47012 38388 47294
rect 39116 47346 39172 48076
rect 40796 48038 40852 48076
rect 39116 47294 39118 47346
rect 39170 47294 39172 47346
rect 39116 47282 39172 47294
rect 38332 46946 38388 46956
rect 41580 47124 41636 47134
rect 37100 46846 37102 46898
rect 37154 46846 37156 46898
rect 37100 46834 37156 46846
rect 32732 46498 32788 46508
rect 38332 46786 38388 46798
rect 38332 46734 38334 46786
rect 38386 46734 38388 46786
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 38332 46002 38388 46734
rect 41580 46674 41636 47068
rect 41692 47012 41748 47022
rect 41692 46786 41748 46956
rect 41692 46734 41694 46786
rect 41746 46734 41748 46786
rect 41692 46722 41748 46734
rect 42028 46786 42084 46798
rect 42028 46734 42030 46786
rect 42082 46734 42084 46786
rect 41580 46622 41582 46674
rect 41634 46622 41636 46674
rect 41580 46610 41636 46622
rect 40796 46562 40852 46574
rect 40796 46510 40798 46562
rect 40850 46510 40852 46562
rect 38332 45950 38334 46002
rect 38386 45950 38388 46002
rect 38332 45938 38388 45950
rect 40460 46002 40516 46014
rect 40460 45950 40462 46002
rect 40514 45950 40516 46002
rect 33628 45890 33684 45902
rect 33628 45838 33630 45890
rect 33682 45838 33684 45890
rect 32956 45778 33012 45790
rect 32956 45726 32958 45778
rect 33010 45726 33012 45778
rect 32956 45668 33012 45726
rect 32956 45602 33012 45612
rect 33628 45668 33684 45838
rect 37660 45892 37716 45902
rect 37660 45798 37716 45836
rect 34188 45668 34244 45678
rect 33628 45666 34244 45668
rect 33628 45614 34190 45666
rect 34242 45614 34244 45666
rect 33628 45612 34244 45614
rect 31724 45378 31780 45388
rect 31276 45054 31278 45106
rect 31330 45054 31332 45106
rect 31276 45042 31332 45054
rect 31164 43710 31166 43762
rect 31218 43710 31220 43762
rect 31164 43698 31220 43710
rect 30716 43374 30718 43426
rect 30770 43374 30772 43426
rect 30716 43362 30772 43374
rect 27804 42130 27860 42140
rect 33628 42754 33684 45612
rect 34188 45602 34244 45612
rect 35308 45108 35364 45118
rect 40460 45108 40516 45950
rect 40796 45892 40852 46510
rect 40796 45826 40852 45836
rect 41020 45892 41076 45902
rect 41020 45798 41076 45836
rect 41468 45892 41524 45902
rect 40796 45332 40852 45342
rect 40796 45238 40852 45276
rect 35308 45106 35588 45108
rect 35308 45054 35310 45106
rect 35362 45054 35588 45106
rect 35308 45052 35588 45054
rect 35308 45042 35364 45052
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 33964 44100 34020 44110
rect 33964 44098 34468 44100
rect 33964 44046 33966 44098
rect 34018 44046 34468 44098
rect 33964 44044 34468 44046
rect 33964 44034 34020 44044
rect 34412 42866 34468 44044
rect 34412 42814 34414 42866
rect 34466 42814 34468 42866
rect 34412 42802 34468 42814
rect 35084 43538 35140 43550
rect 35084 43486 35086 43538
rect 35138 43486 35140 43538
rect 33628 42702 33630 42754
rect 33682 42702 33684 42754
rect 31612 42084 31668 42094
rect 32620 42084 32676 42094
rect 29260 41972 29316 41982
rect 27300 40348 27412 40404
rect 28588 40516 28644 40526
rect 27244 40310 27300 40348
rect 27132 40124 27860 40180
rect 26908 39006 26910 39058
rect 26962 39006 26964 39058
rect 26908 38994 26964 39006
rect 27020 39732 27076 39742
rect 26796 38836 26852 38846
rect 26796 38742 26852 38780
rect 27020 38834 27076 39676
rect 27804 39730 27860 40124
rect 27804 39678 27806 39730
rect 27858 39678 27860 39730
rect 27804 39666 27860 39678
rect 27020 38782 27022 38834
rect 27074 38782 27076 38834
rect 27020 38770 27076 38782
rect 27692 39620 27748 39630
rect 27692 38836 27748 39564
rect 28588 39618 28644 40460
rect 29260 40516 29316 41916
rect 29932 41860 29988 41870
rect 29932 41858 30212 41860
rect 29932 41806 29934 41858
rect 29986 41806 30212 41858
rect 29932 41804 30212 41806
rect 29932 41794 29988 41804
rect 30156 41074 30212 41804
rect 31612 41186 31668 42028
rect 32284 42082 32676 42084
rect 32284 42030 32622 42082
rect 32674 42030 32676 42082
rect 32284 42028 32676 42030
rect 32060 41858 32116 41870
rect 32060 41806 32062 41858
rect 32114 41806 32116 41858
rect 32060 41412 32116 41806
rect 32060 41346 32116 41356
rect 32284 41298 32340 42028
rect 32620 42018 32676 42028
rect 33628 42084 33684 42702
rect 32284 41246 32286 41298
rect 32338 41246 32340 41298
rect 32284 41234 32340 41246
rect 31612 41134 31614 41186
rect 31666 41134 31668 41186
rect 31612 41122 31668 41134
rect 30156 41022 30158 41074
rect 30210 41022 30212 41074
rect 30156 41010 30212 41022
rect 29260 40422 29316 40460
rect 33628 40402 33684 42028
rect 34300 42082 34356 42094
rect 34300 42030 34302 42082
rect 34354 42030 34356 42082
rect 34300 40516 34356 42030
rect 34748 42084 34804 42094
rect 34748 41990 34804 42028
rect 34412 41300 34468 41310
rect 34412 41206 34468 41244
rect 34412 40516 34468 40526
rect 34300 40514 34468 40516
rect 34300 40462 34414 40514
rect 34466 40462 34468 40514
rect 34300 40460 34468 40462
rect 34412 40450 34468 40460
rect 33628 40350 33630 40402
rect 33682 40350 33684 40402
rect 33628 40338 33684 40350
rect 31948 39788 32564 39844
rect 28588 39566 28590 39618
rect 28642 39566 28644 39618
rect 28588 39554 28644 39566
rect 29708 39620 29764 39630
rect 29708 39526 29764 39564
rect 30380 39506 30436 39518
rect 30380 39454 30382 39506
rect 30434 39454 30436 39506
rect 27244 38612 27300 38622
rect 27244 38610 27412 38612
rect 27244 38558 27246 38610
rect 27298 38558 27412 38610
rect 27244 38556 27412 38558
rect 27244 38546 27300 38556
rect 24892 37378 24948 37390
rect 24892 37326 24894 37378
rect 24946 37326 24948 37378
rect 24892 36596 24948 37326
rect 26684 37266 26740 37436
rect 26684 37214 26686 37266
rect 26738 37214 26740 37266
rect 26684 37202 26740 37214
rect 24892 36530 24948 36540
rect 25340 36596 25396 36606
rect 27356 36596 27412 38556
rect 27468 38610 27524 38622
rect 27468 38558 27470 38610
rect 27522 38558 27524 38610
rect 27468 38162 27524 38558
rect 27468 38110 27470 38162
rect 27522 38110 27524 38162
rect 27468 38098 27524 38110
rect 27692 37380 27748 38780
rect 28364 38836 28420 38846
rect 28364 38742 28420 38780
rect 29036 38722 29092 38734
rect 29036 38670 29038 38722
rect 29090 38670 29092 38722
rect 29036 38668 29092 38670
rect 29036 38612 29652 38668
rect 29596 37938 29652 38612
rect 29596 37886 29598 37938
rect 29650 37886 29652 37938
rect 29596 37874 29652 37886
rect 30380 37938 30436 39454
rect 31612 38836 31668 38846
rect 31612 38742 31668 38780
rect 31164 38722 31220 38734
rect 31164 38670 31166 38722
rect 31218 38670 31220 38722
rect 31164 38668 31220 38670
rect 31164 38612 31556 38668
rect 30380 37886 30382 37938
rect 30434 37886 30436 37938
rect 30380 37874 30436 37886
rect 27916 37826 27972 37838
rect 27916 37774 27918 37826
rect 27970 37774 27972 37826
rect 27916 37380 27972 37774
rect 27692 37378 27972 37380
rect 27692 37326 27694 37378
rect 27746 37326 27972 37378
rect 27692 37324 27972 37326
rect 27692 37314 27748 37324
rect 27468 36596 27524 36606
rect 27356 36594 27524 36596
rect 27356 36542 27470 36594
rect 27522 36542 27524 36594
rect 27356 36540 27524 36542
rect 25340 36502 25396 36540
rect 27468 36530 27524 36540
rect 27916 36594 27972 37324
rect 31500 37268 31556 38612
rect 31724 37268 31780 37278
rect 31500 37266 31780 37268
rect 31500 37214 31726 37266
rect 31778 37214 31780 37266
rect 31500 37212 31780 37214
rect 31724 37202 31780 37212
rect 31948 37266 32004 39788
rect 32508 39730 32564 39788
rect 32508 39678 32510 39730
rect 32562 39678 32564 39730
rect 32508 39666 32564 39678
rect 31948 37214 31950 37266
rect 32002 37214 32004 37266
rect 31948 37202 32004 37214
rect 32172 39620 32228 39630
rect 32172 38050 32228 39564
rect 32956 39620 33012 39630
rect 32956 39526 33012 39564
rect 32844 38948 32900 38958
rect 32844 38162 32900 38892
rect 33628 38948 33684 38958
rect 33628 38854 33684 38892
rect 35084 38836 35140 43486
rect 35532 43428 35588 45052
rect 40460 45042 40516 45052
rect 35980 44996 36036 45006
rect 38108 44996 38164 45006
rect 35980 44994 36260 44996
rect 35980 44942 35982 44994
rect 36034 44942 36260 44994
rect 35980 44940 36260 44942
rect 35980 44930 36036 44940
rect 36204 44210 36260 44940
rect 38108 44902 38164 44940
rect 38556 44994 38612 45006
rect 38556 44942 38558 44994
rect 38610 44942 38612 44994
rect 36204 44158 36206 44210
rect 36258 44158 36260 44210
rect 36204 44146 36260 44158
rect 35756 43428 35812 43438
rect 35532 43426 35812 43428
rect 35532 43374 35758 43426
rect 35810 43374 35812 43426
rect 35532 43372 35812 43374
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35756 42084 35812 43372
rect 36540 42868 36596 42878
rect 35756 42018 35812 42028
rect 35868 42866 36596 42868
rect 35868 42814 36542 42866
rect 36594 42814 36596 42866
rect 35868 42812 36596 42814
rect 35868 41860 35924 42812
rect 36540 42802 36596 42812
rect 37548 42532 37604 42542
rect 37212 42530 37604 42532
rect 37212 42478 37550 42530
rect 37602 42478 37604 42530
rect 37212 42476 37604 42478
rect 36988 42084 37044 42094
rect 36540 41972 36596 41982
rect 36540 41878 36596 41916
rect 35532 41804 35924 41860
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 41412 35252 41422
rect 35196 41318 35252 41356
rect 35532 41410 35588 41804
rect 35532 41358 35534 41410
rect 35586 41358 35588 41410
rect 35532 41346 35588 41358
rect 35308 41300 35364 41310
rect 35308 41206 35364 41244
rect 35756 41188 35812 41198
rect 35756 41186 36596 41188
rect 35756 41134 35758 41186
rect 35810 41134 36596 41186
rect 35756 41132 36596 41134
rect 35756 41122 35812 41132
rect 35644 40962 35700 40974
rect 35644 40910 35646 40962
rect 35698 40910 35700 40962
rect 35644 40292 35700 40910
rect 35644 40226 35700 40236
rect 36540 40290 36596 41132
rect 36988 40626 37044 42028
rect 37212 42082 37268 42476
rect 37548 42466 37604 42476
rect 38108 42532 38164 42542
rect 38556 42532 38612 44942
rect 39676 43652 39732 43662
rect 39452 43650 39732 43652
rect 39452 43598 39678 43650
rect 39730 43598 39732 43650
rect 39452 43596 39732 43598
rect 39452 42866 39508 43596
rect 39676 43586 39732 43596
rect 40236 43540 40292 43550
rect 40236 43428 40292 43484
rect 39452 42814 39454 42866
rect 39506 42814 39508 42866
rect 39452 42802 39508 42814
rect 40012 43426 40292 43428
rect 40012 43374 40238 43426
rect 40290 43374 40292 43426
rect 40012 43372 40292 43374
rect 38108 42530 38612 42532
rect 38108 42478 38110 42530
rect 38162 42478 38612 42530
rect 38108 42476 38612 42478
rect 38780 42754 38836 42766
rect 38780 42702 38782 42754
rect 38834 42702 38836 42754
rect 37212 42030 37214 42082
rect 37266 42030 37268 42082
rect 37212 42018 37268 42030
rect 38108 42084 38164 42476
rect 38108 42018 38164 42028
rect 38780 41972 38836 42702
rect 38108 40964 38164 40974
rect 38108 40962 38612 40964
rect 38108 40910 38110 40962
rect 38162 40910 38612 40962
rect 38108 40908 38612 40910
rect 38108 40898 38164 40908
rect 36988 40574 36990 40626
rect 37042 40574 37044 40626
rect 36988 40562 37044 40574
rect 38556 40514 38612 40908
rect 38556 40462 38558 40514
rect 38610 40462 38612 40514
rect 38556 40450 38612 40462
rect 37884 40404 37940 40414
rect 37884 40310 37940 40348
rect 38780 40404 38836 41916
rect 39340 42084 39396 42094
rect 39340 41858 39396 42028
rect 39340 41806 39342 41858
rect 39394 41806 39396 41858
rect 39340 41794 39396 41806
rect 38780 40338 38836 40348
rect 36540 40238 36542 40290
rect 36594 40238 36596 40290
rect 36540 40226 36596 40238
rect 37324 40292 37380 40302
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35084 38704 35140 38780
rect 36988 38724 37044 38800
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 32844 38110 32846 38162
rect 32898 38110 32900 38162
rect 32844 38098 32900 38110
rect 34972 38164 35028 38174
rect 34972 38070 35028 38108
rect 36316 38164 36372 38174
rect 36316 38070 36372 38108
rect 36652 38164 36708 38174
rect 36652 38070 36708 38108
rect 32172 37998 32174 38050
rect 32226 37998 32228 38050
rect 32172 37268 32228 37998
rect 36428 38052 36484 38062
rect 36428 38050 36596 38052
rect 36428 37998 36430 38050
rect 36482 37998 36596 38050
rect 36428 37996 36596 37998
rect 36428 37986 36484 37996
rect 35532 37826 35588 37838
rect 35532 37774 35534 37826
rect 35586 37774 35588 37826
rect 34636 37380 34692 37390
rect 34636 37286 34692 37324
rect 35532 37380 35588 37774
rect 36540 37604 36596 37996
rect 36764 37940 36820 37950
rect 36764 37846 36820 37884
rect 36540 37548 36820 37604
rect 35532 37314 35588 37324
rect 32172 37202 32228 37212
rect 33852 37268 33908 37278
rect 33852 37174 33908 37212
rect 35084 37268 35140 37278
rect 32508 37156 32564 37166
rect 32508 37062 32564 37100
rect 27916 36542 27918 36594
rect 27970 36542 27972 36594
rect 23548 35634 23604 35644
rect 23772 36482 24612 36484
rect 23772 36430 24558 36482
rect 24610 36430 24612 36482
rect 23772 36428 24612 36430
rect 23100 35138 23380 35140
rect 23100 35086 23102 35138
rect 23154 35086 23380 35138
rect 23100 35084 23380 35086
rect 23100 35074 23156 35084
rect 22540 34914 22596 34926
rect 22764 34916 22820 34926
rect 22540 34862 22542 34914
rect 22594 34862 22596 34914
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 22540 34356 22596 34862
rect 22428 34300 22596 34356
rect 22652 34914 22820 34916
rect 22652 34862 22766 34914
rect 22818 34862 22820 34914
rect 22652 34860 22820 34862
rect 18620 33406 18622 33458
rect 18674 33406 18676 33458
rect 18620 33394 18676 33406
rect 18732 34132 18788 34142
rect 17164 33294 17166 33346
rect 17218 33294 17220 33346
rect 16156 32788 16212 32798
rect 16156 32694 16212 32732
rect 17164 32788 17220 33294
rect 15708 32452 15764 32462
rect 15708 32450 15876 32452
rect 15708 32398 15710 32450
rect 15762 32398 15876 32450
rect 15708 32396 15876 32398
rect 15708 32386 15764 32396
rect 15820 31948 15876 32396
rect 17164 31948 17220 32732
rect 17836 33346 17892 33358
rect 17836 33294 17838 33346
rect 17890 33294 17892 33346
rect 17836 32562 17892 33294
rect 17836 32510 17838 32562
rect 17890 32510 17892 32562
rect 17836 31948 17892 32510
rect 18508 32450 18564 32462
rect 18508 32398 18510 32450
rect 18562 32398 18564 32450
rect 18508 31948 18564 32398
rect 15708 31892 15764 31902
rect 15820 31892 15988 31948
rect 16604 31892 16660 31902
rect 15708 30994 15764 31836
rect 15708 30942 15710 30994
rect 15762 30942 15764 30994
rect 15708 30930 15764 30942
rect 15932 30994 15988 31892
rect 15932 30942 15934 30994
rect 15986 30942 15988 30994
rect 15932 30930 15988 30942
rect 16156 31890 16660 31892
rect 16156 31838 16606 31890
rect 16658 31838 16660 31890
rect 16156 31836 16660 31838
rect 16156 30994 16212 31836
rect 16604 31826 16660 31836
rect 17164 31890 17332 31948
rect 17836 31892 18004 31948
rect 17164 31838 17166 31890
rect 17218 31838 17332 31890
rect 17164 31836 17332 31838
rect 17164 31826 17220 31836
rect 17948 31826 18004 31836
rect 18284 31892 18564 31948
rect 18284 31666 18340 31892
rect 18284 31614 18286 31666
rect 18338 31614 18340 31666
rect 18284 31602 18340 31614
rect 16156 30942 16158 30994
rect 16210 30942 16212 30994
rect 16156 30930 16212 30942
rect 16268 31220 16324 31230
rect 16268 30994 16324 31164
rect 16268 30942 16270 30994
rect 16322 30942 16324 30994
rect 16268 30930 16324 30942
rect 18508 30996 18564 31006
rect 18508 30902 18564 30940
rect 15372 28588 15540 28644
rect 15596 30770 15652 30782
rect 15596 30718 15598 30770
rect 15650 30718 15652 30770
rect 13804 28418 13860 28430
rect 13804 28366 13806 28418
rect 13858 28366 13860 28418
rect 13692 27972 13748 27982
rect 13804 27972 13860 28366
rect 15148 28420 15204 28430
rect 15148 28326 15204 28364
rect 15260 28418 15316 28430
rect 15260 28366 15262 28418
rect 15314 28366 15316 28418
rect 13692 27970 13860 27972
rect 13692 27918 13694 27970
rect 13746 27918 13860 27970
rect 13692 27916 13860 27918
rect 13692 27906 13748 27916
rect 12908 27346 12964 27356
rect 13020 27858 13076 27870
rect 13020 27806 13022 27858
rect 13074 27806 13076 27858
rect 8204 26798 8206 26850
rect 8258 26798 8260 26850
rect 7532 26238 7534 26290
rect 7586 26238 7588 26290
rect 7532 26180 7588 26238
rect 7532 26114 7588 26124
rect 7980 26404 8036 26414
rect 7868 26068 7924 26078
rect 7868 25974 7924 26012
rect 7868 25620 7924 25630
rect 7980 25620 8036 26348
rect 8204 25732 8260 26798
rect 8540 27186 9492 27188
rect 8540 27134 8990 27186
rect 9042 27134 9438 27186
rect 9490 27134 9492 27186
rect 8540 27132 9492 27134
rect 8540 27074 8596 27132
rect 8988 27122 9044 27132
rect 9436 27122 9492 27132
rect 10780 27188 10836 27198
rect 12908 27188 12964 27198
rect 10780 27186 11508 27188
rect 10780 27134 10782 27186
rect 10834 27134 11508 27186
rect 10780 27132 11508 27134
rect 10780 27122 10836 27132
rect 8540 27022 8542 27074
rect 8594 27022 8596 27074
rect 8540 26290 8596 27022
rect 10108 27074 10164 27086
rect 10108 27022 10110 27074
rect 10162 27022 10164 27074
rect 10108 26964 10164 27022
rect 10108 26898 10164 26908
rect 11228 26964 11284 26974
rect 8540 26238 8542 26290
rect 8594 26238 8596 26290
rect 8540 26226 8596 26238
rect 8876 26514 8932 26526
rect 8876 26462 8878 26514
rect 8930 26462 8932 26514
rect 8764 26068 8820 26078
rect 8764 25974 8820 26012
rect 8876 25844 8932 26462
rect 9996 26404 10052 26414
rect 9996 26310 10052 26348
rect 8988 26292 9044 26302
rect 9884 26292 9940 26302
rect 8988 26290 9940 26292
rect 8988 26238 8990 26290
rect 9042 26238 9886 26290
rect 9938 26238 9940 26290
rect 8988 26236 9940 26238
rect 8988 26226 9044 26236
rect 9884 26226 9940 26236
rect 9772 26068 9828 26078
rect 9772 25974 9828 26012
rect 8876 25788 10052 25844
rect 8204 25666 8260 25676
rect 7868 25618 8036 25620
rect 7868 25566 7870 25618
rect 7922 25566 8036 25618
rect 7868 25564 8036 25566
rect 9996 25618 10052 25788
rect 11228 25620 11284 26908
rect 11452 26514 11508 27132
rect 12908 27094 12964 27132
rect 13020 26964 13076 27806
rect 14924 27748 14980 27758
rect 14700 27412 14756 27422
rect 14700 27298 14756 27356
rect 14700 27246 14702 27298
rect 14754 27246 14756 27298
rect 14700 27234 14756 27246
rect 14812 27188 14868 27198
rect 14812 27094 14868 27132
rect 13020 26898 13076 26908
rect 13580 26964 13636 26974
rect 11452 26462 11454 26514
rect 11506 26462 11508 26514
rect 11452 26450 11508 26462
rect 9996 25566 9998 25618
rect 10050 25566 10052 25618
rect 7868 25554 7924 25564
rect 9996 25554 10052 25566
rect 10780 25618 11284 25620
rect 10780 25566 11230 25618
rect 11282 25566 11284 25618
rect 10780 25564 11284 25566
rect 10780 25506 10836 25564
rect 11228 25554 11284 25564
rect 10780 25454 10782 25506
rect 10834 25454 10836 25506
rect 10780 25442 10836 25454
rect 7308 24670 7310 24722
rect 7362 24670 7364 24722
rect 7308 24658 7364 24670
rect 13020 24722 13076 24734
rect 13020 24670 13022 24722
rect 13074 24670 13076 24722
rect 7084 24610 7140 24622
rect 7084 24558 7086 24610
rect 7138 24558 7140 24610
rect 7084 23604 7140 24558
rect 12236 24052 12292 24062
rect 13020 24052 13076 24670
rect 12236 24050 12628 24052
rect 12236 23998 12238 24050
rect 12290 23998 12628 24050
rect 12236 23996 12628 23998
rect 12236 23986 12292 23996
rect 7084 23538 7140 23548
rect 9436 23938 9492 23950
rect 9436 23886 9438 23938
rect 9490 23886 9492 23938
rect 6860 23202 6916 23212
rect 8428 23268 8484 23278
rect 5740 23154 6132 23156
rect 5740 23102 6078 23154
rect 6130 23102 6132 23154
rect 5740 23100 6132 23102
rect 5516 23042 5572 23054
rect 5516 22990 5518 23042
rect 5570 22990 5572 23042
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 5516 22596 5572 22990
rect 5516 22540 5796 22596
rect 3948 22430 3950 22482
rect 4002 22430 4004 22482
rect 3948 22418 4004 22430
rect 2716 21858 2772 21868
rect 4732 22370 4788 22382
rect 4732 22318 4734 22370
rect 4786 22318 4788 22370
rect 4732 21924 4788 22318
rect 4732 21858 4788 21868
rect 4956 21924 5012 21934
rect 4956 21810 5012 21868
rect 4956 21758 4958 21810
rect 5010 21758 5012 21810
rect 4956 21746 5012 21758
rect 5628 21924 5684 21934
rect 2492 21588 2548 21598
rect 2492 21474 2548 21532
rect 2492 21422 2494 21474
rect 2546 21422 2548 21474
rect 2492 21410 2548 21422
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 5628 20914 5684 21868
rect 5628 20862 5630 20914
rect 5682 20862 5684 20914
rect 2156 20132 2324 20188
rect 2828 20580 2884 20590
rect 2156 20018 2212 20132
rect 2156 19966 2158 20018
rect 2210 19966 2212 20018
rect 2156 19234 2212 19966
rect 2828 19346 2884 20524
rect 3164 20578 3220 20590
rect 3164 20526 3166 20578
rect 3218 20526 3220 20578
rect 3164 20188 3220 20526
rect 3836 20580 3892 20590
rect 3836 20486 3892 20524
rect 2940 20132 3220 20188
rect 2940 20130 2996 20132
rect 2940 20078 2942 20130
rect 2994 20078 2996 20130
rect 2940 20066 2996 20078
rect 5628 20018 5684 20862
rect 5740 20188 5796 22540
rect 6076 21924 6132 23100
rect 6636 23044 6692 23054
rect 6636 22370 6692 22988
rect 6860 23044 6916 23054
rect 6860 23042 7364 23044
rect 6860 22990 6862 23042
rect 6914 22990 7364 23042
rect 6860 22988 7364 22990
rect 6860 22978 6916 22988
rect 6636 22318 6638 22370
rect 6690 22318 6692 22370
rect 6636 22306 6692 22318
rect 6076 21858 6132 21868
rect 7308 21810 7364 22988
rect 8428 22484 8484 23212
rect 8988 23044 9044 23054
rect 8988 23042 9156 23044
rect 8988 22990 8990 23042
rect 9042 22990 9156 23042
rect 8988 22988 9156 22990
rect 8988 22978 9044 22988
rect 8428 22352 8484 22428
rect 8988 22484 9044 22494
rect 7308 21758 7310 21810
rect 7362 21758 7364 21810
rect 7308 21746 7364 21758
rect 6524 20578 6580 20590
rect 6524 20526 6526 20578
rect 6578 20526 6580 20578
rect 5740 20132 6244 20188
rect 5628 19966 5630 20018
rect 5682 19966 5684 20018
rect 5068 19906 5124 19918
rect 5068 19854 5070 19906
rect 5122 19854 5124 19906
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 5068 19460 5124 19854
rect 5068 19394 5124 19404
rect 2828 19294 2830 19346
rect 2882 19294 2884 19346
rect 2828 19282 2884 19294
rect 4956 19348 5012 19358
rect 4956 19254 5012 19292
rect 2156 19182 2158 19234
rect 2210 19182 2212 19234
rect 2156 19170 2212 19182
rect 5292 18676 5348 18686
rect 5628 18676 5684 19966
rect 6188 19684 6244 20132
rect 6412 20132 6468 20142
rect 6524 20132 6580 20526
rect 6412 20130 6580 20132
rect 6412 20078 6414 20130
rect 6466 20078 6580 20130
rect 6412 20076 6580 20078
rect 8988 20130 9044 22428
rect 9100 22372 9156 22988
rect 9100 22306 9156 22316
rect 9436 21588 9492 23886
rect 10108 23828 10164 23838
rect 10108 23826 10388 23828
rect 10108 23774 10110 23826
rect 10162 23774 10388 23826
rect 10108 23772 10388 23774
rect 10108 23762 10164 23772
rect 10332 23378 10388 23772
rect 10332 23326 10334 23378
rect 10386 23326 10388 23378
rect 10332 23314 10388 23326
rect 11228 23380 11284 23390
rect 9660 23268 9716 23278
rect 9660 23174 9716 23212
rect 11228 23044 11284 23324
rect 11228 22978 11284 22988
rect 11788 23380 11844 23390
rect 9436 21522 9492 21532
rect 9884 21588 9940 21598
rect 9884 21494 9940 21532
rect 10556 21474 10612 21486
rect 10556 21422 10558 21474
rect 10610 21422 10612 21474
rect 9100 20804 9156 20814
rect 9100 20802 9716 20804
rect 9100 20750 9102 20802
rect 9154 20750 9716 20802
rect 9100 20748 9716 20750
rect 9100 20738 9156 20748
rect 8988 20078 8990 20130
rect 9042 20078 9044 20130
rect 6412 20066 6468 20076
rect 8988 20066 9044 20078
rect 8540 19906 8596 19918
rect 8540 19854 8542 19906
rect 8594 19854 8596 19906
rect 6188 19628 6580 19684
rect 6300 19460 6356 19470
rect 6300 19366 6356 19404
rect 6524 19458 6580 19628
rect 6524 19406 6526 19458
rect 6578 19406 6580 19458
rect 6524 19394 6580 19406
rect 6748 19460 6804 19470
rect 6748 19366 6804 19404
rect 8540 19460 8596 19854
rect 8540 19394 8596 19404
rect 6076 19348 6132 19358
rect 6076 19254 6132 19292
rect 9660 19234 9716 20748
rect 9772 20690 9828 20702
rect 9772 20638 9774 20690
rect 9826 20638 9828 20690
rect 9772 20244 9828 20638
rect 9884 20244 9940 20254
rect 9772 20242 9940 20244
rect 9772 20190 9886 20242
rect 9938 20190 9940 20242
rect 9772 20188 9940 20190
rect 10556 20244 10612 21422
rect 10668 20244 10724 20254
rect 10556 20242 10724 20244
rect 10556 20190 10670 20242
rect 10722 20190 10724 20242
rect 10556 20188 10724 20190
rect 9884 20178 9940 20188
rect 10668 20178 10724 20188
rect 9660 19182 9662 19234
rect 9714 19182 9716 19234
rect 5292 18674 5684 18676
rect 5292 18622 5294 18674
rect 5346 18622 5684 18674
rect 5292 18620 5684 18622
rect 7196 19010 7252 19022
rect 7196 18958 7198 19010
rect 7250 18958 7252 19010
rect 5292 18610 5348 18620
rect 2156 18452 2212 18462
rect 7196 18452 7252 18958
rect 7644 18452 7700 18462
rect 7196 18450 7700 18452
rect 7196 18398 7646 18450
rect 7698 18398 7700 18450
rect 7196 18396 7700 18398
rect 2156 16770 2212 18396
rect 7644 18386 7700 18396
rect 7868 18452 7924 18462
rect 7868 18358 7924 18396
rect 8204 18452 8260 18462
rect 8204 18450 8596 18452
rect 8204 18398 8206 18450
rect 8258 18398 8596 18450
rect 8204 18396 8596 18398
rect 8204 18386 8260 18396
rect 8428 18226 8484 18238
rect 8428 18174 8430 18226
rect 8482 18174 8484 18226
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 8316 17668 8372 17678
rect 6524 17442 6580 17454
rect 6524 17390 6526 17442
rect 6578 17390 6580 17442
rect 6412 16996 6468 17006
rect 6524 16996 6580 17390
rect 6412 16994 6580 16996
rect 6412 16942 6414 16994
rect 6466 16942 6580 16994
rect 6412 16940 6580 16942
rect 6412 16930 6468 16940
rect 5068 16882 5124 16894
rect 5068 16830 5070 16882
rect 5122 16830 5124 16882
rect 2156 16718 2158 16770
rect 2210 16718 2212 16770
rect 2156 16706 2212 16718
rect 4284 16770 4340 16782
rect 4284 16718 4286 16770
rect 4338 16718 4340 16770
rect 4284 15988 4340 16718
rect 5068 16772 5124 16830
rect 5068 16706 5124 16716
rect 5740 16882 5796 16894
rect 5740 16830 5742 16882
rect 5794 16830 5796 16882
rect 5740 16772 5796 16830
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 5628 16212 5684 16222
rect 5740 16212 5796 16716
rect 5628 16210 5796 16212
rect 5628 16158 5630 16210
rect 5682 16158 5796 16210
rect 5628 16156 5796 16158
rect 5628 16146 5684 16156
rect 4508 15988 4564 15998
rect 4284 15986 4564 15988
rect 4284 15934 4510 15986
rect 4562 15934 4564 15986
rect 4284 15932 4564 15934
rect 4508 15922 4564 15932
rect 7980 15092 8036 15102
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 7980 14530 8036 15036
rect 7980 14478 7982 14530
rect 8034 14478 8036 14530
rect 7980 14466 8036 14478
rect 6972 13860 7028 13870
rect 8092 13860 8148 13870
rect 6972 13858 8148 13860
rect 6972 13806 6974 13858
rect 7026 13806 8094 13858
rect 8146 13806 8148 13858
rect 6972 13804 8148 13806
rect 6972 13794 7028 13804
rect 3500 13746 3556 13758
rect 3500 13694 3502 13746
rect 3554 13694 3556 13746
rect 1932 12068 1988 12078
rect 1932 9826 1988 12012
rect 3500 12068 3556 13694
rect 4172 13634 4228 13646
rect 4172 13582 4174 13634
rect 4226 13582 4228 13634
rect 4172 13076 4228 13582
rect 6300 13636 6356 13646
rect 6300 13542 6356 13580
rect 6860 13636 6916 13646
rect 6860 13542 6916 13580
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4172 13010 4228 13020
rect 6972 13076 7028 13086
rect 6972 12982 7028 13020
rect 6076 12964 6132 12974
rect 6076 12870 6132 12908
rect 7084 12962 7140 13804
rect 8092 13794 8148 13804
rect 7756 13634 7812 13646
rect 7756 13582 7758 13634
rect 7810 13582 7812 13634
rect 7084 12910 7086 12962
rect 7138 12910 7140 12962
rect 7084 12898 7140 12910
rect 7308 12964 7364 12974
rect 6636 12850 6692 12862
rect 6636 12798 6638 12850
rect 6690 12798 6692 12850
rect 4284 12740 4340 12750
rect 3500 12002 3556 12012
rect 3948 12068 4004 12078
rect 3948 11974 4004 12012
rect 2828 10610 2884 10622
rect 2828 10558 2830 10610
rect 2882 10558 2884 10610
rect 2828 10500 2884 10558
rect 3164 10612 3220 10622
rect 2828 10164 2884 10444
rect 1932 9774 1934 9826
rect 1986 9774 1988 9826
rect 1932 9762 1988 9774
rect 2492 10108 2884 10164
rect 3052 10498 3108 10510
rect 3052 10446 3054 10498
rect 3106 10446 3108 10498
rect 2156 8258 2212 8270
rect 2156 8206 2158 8258
rect 2210 8206 2212 8258
rect 2156 7588 2212 8206
rect 2156 7522 2212 7532
rect 2492 7476 2548 10108
rect 3052 10052 3108 10446
rect 2604 9996 3108 10052
rect 2604 9938 2660 9996
rect 3164 9940 3220 10556
rect 3388 10610 3444 10622
rect 3388 10558 3390 10610
rect 3442 10558 3444 10610
rect 3388 10388 3444 10558
rect 4284 10612 4340 12684
rect 5740 12740 5796 12750
rect 5740 12646 5796 12684
rect 6636 12740 6692 12798
rect 6636 12674 6692 12684
rect 6860 12852 6916 12862
rect 6860 12738 6916 12796
rect 6860 12686 6862 12738
rect 6914 12686 6916 12738
rect 6860 12292 6916 12686
rect 7196 12738 7252 12750
rect 7196 12686 7198 12738
rect 7250 12686 7252 12738
rect 7196 12404 7252 12686
rect 7196 12338 7252 12348
rect 6636 12236 6916 12292
rect 5740 12068 5796 12078
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 5740 11394 5796 12012
rect 5740 11342 5742 11394
rect 5794 11342 5796 11394
rect 5740 11330 5796 11342
rect 6524 11284 6580 11294
rect 6524 11190 6580 11228
rect 4396 10612 4452 10622
rect 4284 10556 4396 10612
rect 4396 10518 4452 10556
rect 6636 10610 6692 12236
rect 6748 11284 6804 11294
rect 6748 10834 6804 11228
rect 6748 10782 6750 10834
rect 6802 10782 6804 10834
rect 6748 10770 6804 10782
rect 6636 10558 6638 10610
rect 6690 10558 6692 10610
rect 6636 10546 6692 10558
rect 6972 10612 7028 10622
rect 7308 10612 7364 12908
rect 7756 12964 7812 13582
rect 7756 12898 7812 12908
rect 8204 12852 8260 12862
rect 7756 12740 7812 12750
rect 7756 12646 7812 12684
rect 8204 11396 8260 12796
rect 8316 12180 8372 17612
rect 8428 13860 8484 18174
rect 8540 16770 8596 18396
rect 8988 16884 9044 16894
rect 8540 16718 8542 16770
rect 8594 16718 8596 16770
rect 8540 16706 8596 16718
rect 8764 16828 8988 16884
rect 8764 16772 8820 16828
rect 8988 16790 9044 16828
rect 9660 16884 9716 19182
rect 10444 19124 10500 19134
rect 10444 19122 10724 19124
rect 10444 19070 10446 19122
rect 10498 19070 10724 19122
rect 10444 19068 10724 19070
rect 10444 19058 10500 19068
rect 10668 18674 10724 19068
rect 10668 18622 10670 18674
rect 10722 18622 10724 18674
rect 10668 18610 10724 18622
rect 11788 17780 11844 23324
rect 12012 23156 12068 23166
rect 12012 23062 12068 23100
rect 12348 22596 12404 22606
rect 11900 22594 12404 22596
rect 11900 22542 12350 22594
rect 12402 22542 12404 22594
rect 11900 22540 12404 22542
rect 11900 20914 11956 22540
rect 12348 22530 12404 22540
rect 12572 22594 12628 23996
rect 12908 23828 12964 23838
rect 12908 23734 12964 23772
rect 13020 23380 13076 23996
rect 13020 23314 13076 23324
rect 13580 23940 13636 26908
rect 14924 26964 14980 27692
rect 15260 27636 15316 28366
rect 15148 27580 15316 27636
rect 15036 27300 15092 27310
rect 15036 27206 15092 27244
rect 13692 25284 13748 25294
rect 13692 25282 13860 25284
rect 13692 25230 13694 25282
rect 13746 25230 13860 25282
rect 13692 25228 13860 25230
rect 13692 25218 13748 25228
rect 13692 23940 13748 23950
rect 13580 23938 13748 23940
rect 13580 23886 13694 23938
rect 13746 23886 13748 23938
rect 13580 23884 13748 23886
rect 13356 23268 13412 23278
rect 13356 23174 13412 23212
rect 12684 23156 12740 23166
rect 12684 23062 12740 23100
rect 13132 23156 13188 23166
rect 12572 22542 12574 22594
rect 12626 22542 12628 22594
rect 12572 22530 12628 22542
rect 12012 22372 12068 22410
rect 12012 22306 12068 22316
rect 12124 22372 12180 22382
rect 12124 22370 12292 22372
rect 12124 22318 12126 22370
rect 12178 22318 12292 22370
rect 12124 22316 12292 22318
rect 12124 22306 12180 22316
rect 12236 21924 12292 22316
rect 12684 22260 12740 22270
rect 12684 22258 12852 22260
rect 12684 22206 12686 22258
rect 12738 22206 12852 22258
rect 12684 22204 12852 22206
rect 12684 22194 12740 22204
rect 12236 21868 12740 21924
rect 12684 21474 12740 21868
rect 12684 21422 12686 21474
rect 12738 21422 12740 21474
rect 12684 21410 12740 21422
rect 11900 20862 11902 20914
rect 11954 20862 11956 20914
rect 11900 20850 11956 20862
rect 12348 20580 12404 20590
rect 12348 20486 12404 20524
rect 12796 20188 12852 22204
rect 13132 21810 13188 23100
rect 13580 23156 13636 23884
rect 13692 23874 13748 23884
rect 13804 23268 13860 25228
rect 14924 24834 14980 26908
rect 15148 26850 15204 27580
rect 15148 26798 15150 26850
rect 15202 26798 15204 26850
rect 15148 26786 15204 26798
rect 15260 27074 15316 27086
rect 15260 27022 15262 27074
rect 15314 27022 15316 27074
rect 14924 24782 14926 24834
rect 14978 24782 14980 24834
rect 14476 23828 14532 23838
rect 14476 23734 14532 23772
rect 13804 23202 13860 23212
rect 14588 23380 14644 23390
rect 13580 22482 13636 23100
rect 13580 22430 13582 22482
rect 13634 22430 13636 22482
rect 13580 22418 13636 22430
rect 14588 22372 14644 23324
rect 14924 23380 14980 24782
rect 14924 23314 14980 23324
rect 15260 23156 15316 27022
rect 15372 23268 15428 28588
rect 15484 28420 15540 28430
rect 15596 28420 15652 30718
rect 16380 30324 16436 30334
rect 16380 30210 16436 30268
rect 16380 30158 16382 30210
rect 16434 30158 16436 30210
rect 16380 30146 16436 30158
rect 16716 30324 16772 30334
rect 16716 28642 16772 30268
rect 18620 30324 18676 30334
rect 17052 30100 17108 30110
rect 17052 30098 17780 30100
rect 17052 30046 17054 30098
rect 17106 30046 17780 30098
rect 17052 30044 17780 30046
rect 17052 30034 17108 30044
rect 17724 29650 17780 30044
rect 17724 29598 17726 29650
rect 17778 29598 17780 29650
rect 17724 29586 17780 29598
rect 16940 29540 16996 29550
rect 16940 29538 17444 29540
rect 16940 29486 16942 29538
rect 16994 29486 17444 29538
rect 16940 29484 17444 29486
rect 16940 29474 16996 29484
rect 17388 28754 17444 29484
rect 18620 29426 18676 30268
rect 18620 29374 18622 29426
rect 18674 29374 18676 29426
rect 18620 29362 18676 29374
rect 17388 28702 17390 28754
rect 17442 28702 17444 28754
rect 17388 28690 17444 28702
rect 18732 28756 18788 34076
rect 19628 34130 19684 34142
rect 19628 34078 19630 34130
rect 19682 34078 19684 34130
rect 19404 31892 19460 31902
rect 19404 31798 19460 31836
rect 19628 31892 19684 34078
rect 20412 34020 20468 34030
rect 20412 34018 21700 34020
rect 20412 33966 20414 34018
rect 20466 33966 21700 34018
rect 20412 33964 21700 33966
rect 20412 33954 20468 33964
rect 20748 33684 20804 33694
rect 20748 33458 20804 33628
rect 20748 33406 20750 33458
rect 20802 33406 20804 33458
rect 20748 33394 20804 33406
rect 21644 33234 21700 33964
rect 22428 33684 22484 34300
rect 22652 34244 22708 34860
rect 22764 34850 22820 34860
rect 22540 34188 22708 34244
rect 22540 34018 22596 34188
rect 22988 34020 23044 34030
rect 22540 33966 22542 34018
rect 22594 33966 22596 34018
rect 22540 33954 22596 33966
rect 22652 34018 23044 34020
rect 22652 33966 22990 34018
rect 23042 33966 23044 34018
rect 22652 33964 23044 33966
rect 22428 33618 22484 33628
rect 21644 33182 21646 33234
rect 21698 33182 21700 33234
rect 21644 33170 21700 33182
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 21084 32564 21140 32574
rect 22092 32564 22148 32574
rect 22652 32564 22708 33964
rect 22988 33954 23044 33964
rect 23772 33346 23828 36428
rect 24556 36418 24612 36428
rect 24444 35700 24500 35710
rect 24444 35606 24500 35644
rect 27916 35700 27972 36542
rect 31500 37044 31556 37054
rect 29596 36260 29652 36270
rect 29372 36258 29652 36260
rect 29372 36206 29598 36258
rect 29650 36206 29652 36258
rect 29372 36204 29652 36206
rect 29372 35810 29428 36204
rect 29596 36194 29652 36204
rect 29372 35758 29374 35810
rect 29426 35758 29428 35810
rect 29372 35746 29428 35758
rect 23996 35588 24052 35598
rect 23996 35494 24052 35532
rect 24668 34692 24724 34702
rect 24444 34690 24724 34692
rect 24444 34638 24670 34690
rect 24722 34638 24724 34690
rect 24444 34636 24724 34638
rect 24444 33458 24500 34636
rect 24668 34626 24724 34636
rect 24444 33406 24446 33458
rect 24498 33406 24500 33458
rect 24444 33394 24500 33406
rect 26572 33458 26628 33470
rect 26572 33406 26574 33458
rect 26626 33406 26628 33458
rect 23772 33294 23774 33346
rect 23826 33294 23828 33346
rect 23772 33282 23828 33294
rect 22988 33124 23044 33134
rect 22764 33122 23044 33124
rect 22764 33070 22990 33122
rect 23042 33070 23044 33122
rect 22764 33068 23044 33070
rect 22764 32674 22820 33068
rect 22988 33058 23044 33068
rect 22764 32622 22766 32674
rect 22818 32622 22820 32674
rect 22764 32610 22820 32622
rect 20860 32562 22708 32564
rect 20860 32510 21086 32562
rect 21138 32510 22094 32562
rect 22146 32510 22708 32562
rect 20860 32508 22708 32510
rect 20636 32452 20692 32462
rect 19628 31826 19684 31836
rect 20524 32450 20692 32452
rect 20524 32398 20638 32450
rect 20690 32398 20692 32450
rect 20524 32396 20692 32398
rect 19292 31556 19348 31566
rect 19068 30996 19124 31006
rect 19068 30902 19124 30940
rect 19180 30436 19236 30446
rect 19180 30322 19236 30380
rect 19180 30270 19182 30322
rect 19234 30270 19236 30322
rect 19180 30258 19236 30270
rect 19292 29538 19348 31500
rect 20300 31556 20356 31566
rect 20300 31462 20356 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20188 30436 20244 30446
rect 20188 30342 20244 30380
rect 20300 30324 20356 30334
rect 20076 30212 20132 30222
rect 20076 30118 20132 30156
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20300 29652 20356 30268
rect 19292 29486 19294 29538
rect 19346 29486 19348 29538
rect 19292 29474 19348 29486
rect 20076 29596 20356 29652
rect 20412 30210 20468 30222
rect 20412 30158 20414 30210
rect 20466 30158 20468 30210
rect 18732 28690 18788 28700
rect 19516 28754 19572 28766
rect 19516 28702 19518 28754
rect 19570 28702 19572 28754
rect 16716 28590 16718 28642
rect 16770 28590 16772 28642
rect 16716 28578 16772 28590
rect 15484 28418 15652 28420
rect 15484 28366 15486 28418
rect 15538 28366 15652 28418
rect 15484 28364 15652 28366
rect 15708 28530 15764 28542
rect 15708 28478 15710 28530
rect 15762 28478 15764 28530
rect 15484 28354 15540 28364
rect 15708 28084 15764 28478
rect 19516 28532 19572 28702
rect 20076 28754 20132 29596
rect 20076 28702 20078 28754
rect 20130 28702 20132 28754
rect 20076 28690 20132 28702
rect 19516 28466 19572 28476
rect 20412 28532 20468 30158
rect 20524 30212 20580 32396
rect 20636 32386 20692 32396
rect 20860 31892 20916 32508
rect 21084 32498 21140 32508
rect 20860 31760 20916 31836
rect 21644 31554 21700 32508
rect 22092 32498 22148 32508
rect 24892 32452 24948 32462
rect 24892 32358 24948 32396
rect 26236 32450 26292 32462
rect 26236 32398 26238 32450
rect 26290 32398 26292 32450
rect 21644 31502 21646 31554
rect 21698 31502 21700 31554
rect 21644 31106 21700 31502
rect 21644 31054 21646 31106
rect 21698 31054 21700 31106
rect 20636 30324 20692 30334
rect 21644 30324 21700 31054
rect 24108 31778 24164 31790
rect 24108 31726 24110 31778
rect 24162 31726 24164 31778
rect 20636 30322 21476 30324
rect 20636 30270 20638 30322
rect 20690 30270 21476 30322
rect 20636 30268 21476 30270
rect 20636 30258 20692 30268
rect 20524 30146 20580 30156
rect 20412 28466 20468 28476
rect 20748 30098 20804 30110
rect 20748 30046 20750 30098
rect 20802 30046 20804 30098
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 15708 28018 15764 28028
rect 20748 27858 20804 30046
rect 21420 29314 21476 30268
rect 21700 30268 22036 30324
rect 21644 30192 21700 30268
rect 21980 29428 22036 30268
rect 23324 29988 23380 29998
rect 22764 29986 23380 29988
rect 22764 29934 23326 29986
rect 23378 29934 23380 29986
rect 22764 29932 23380 29934
rect 22764 29538 22820 29932
rect 23324 29922 23380 29932
rect 22764 29486 22766 29538
rect 22818 29486 22820 29538
rect 22764 29474 22820 29486
rect 21420 29262 21422 29314
rect 21474 29262 21476 29314
rect 21420 29250 21476 29262
rect 21756 29426 22036 29428
rect 21756 29374 21982 29426
rect 22034 29374 22036 29426
rect 21756 29372 22036 29374
rect 21756 28754 21812 29372
rect 21980 29362 22036 29372
rect 24108 29428 24164 31726
rect 24780 31666 24836 31678
rect 24780 31614 24782 31666
rect 24834 31614 24836 31666
rect 24780 30098 24836 31614
rect 26236 30996 26292 32398
rect 26572 31948 26628 33406
rect 27804 33460 27860 33470
rect 27916 33460 27972 35644
rect 28588 35700 28644 35710
rect 28588 35606 28644 35644
rect 31500 35586 31556 36988
rect 32172 37044 32228 37054
rect 32396 37044 32452 37054
rect 32172 36950 32228 36988
rect 32284 37042 32452 37044
rect 32284 36990 32398 37042
rect 32450 36990 32452 37042
rect 32284 36988 32452 36990
rect 31948 35700 32004 35710
rect 31948 35606 32004 35644
rect 31500 35534 31502 35586
rect 31554 35534 31556 35586
rect 31500 35522 31556 35534
rect 30156 34690 30212 34702
rect 30156 34638 30158 34690
rect 30210 34638 30212 34690
rect 30044 34244 30100 34254
rect 30156 34244 30212 34638
rect 30044 34242 30212 34244
rect 30044 34190 30046 34242
rect 30098 34190 30212 34242
rect 30044 34188 30212 34190
rect 30044 34178 30100 34188
rect 27804 33458 27972 33460
rect 27804 33406 27806 33458
rect 27858 33406 27972 33458
rect 27804 33404 27972 33406
rect 29372 34130 29428 34142
rect 29372 34078 29374 34130
rect 29426 34078 29428 34130
rect 27804 33394 27860 33404
rect 27244 33124 27300 33134
rect 27244 33122 28420 33124
rect 27244 33070 27246 33122
rect 27298 33070 28420 33122
rect 27244 33068 28420 33070
rect 27244 33058 27300 33068
rect 28364 32674 28420 33068
rect 29372 32788 29428 34078
rect 32172 34020 32228 34030
rect 32284 34020 32340 36988
rect 32396 36978 32452 36988
rect 35084 36708 35140 37212
rect 36764 37154 36820 37548
rect 36764 37102 36766 37154
rect 36818 37102 36820 37154
rect 36764 37090 36820 37102
rect 36988 37268 37044 38668
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35084 36652 35364 36708
rect 35308 36594 35364 36652
rect 35308 36542 35310 36594
rect 35362 36542 35364 36594
rect 35308 36530 35364 36542
rect 36988 36596 37044 37212
rect 37324 37266 37380 40236
rect 37660 39394 37716 39406
rect 37660 39342 37662 39394
rect 37714 39342 37716 39394
rect 37660 38612 37716 39342
rect 40012 39394 40068 43372
rect 40236 43362 40292 43372
rect 40684 42756 40740 42766
rect 40684 40290 40740 42700
rect 41468 41972 41524 45836
rect 41804 45778 41860 45790
rect 41804 45726 41806 45778
rect 41858 45726 41860 45778
rect 41804 45332 41860 45726
rect 42028 45668 42084 46734
rect 42028 45602 42084 45612
rect 41804 45266 41860 45276
rect 42028 45444 42084 45454
rect 41580 45108 41636 45118
rect 41580 45014 41636 45052
rect 42028 45106 42084 45388
rect 42028 45054 42030 45106
rect 42082 45054 42084 45106
rect 42028 45042 42084 45054
rect 41804 44996 41860 45006
rect 41804 44902 41860 44940
rect 42140 43540 42196 49756
rect 42252 49718 42308 49756
rect 42476 48132 42532 48142
rect 42364 46676 42420 46686
rect 42364 46582 42420 46620
rect 42364 45668 42420 45678
rect 42364 45218 42420 45612
rect 42364 45166 42366 45218
rect 42418 45166 42420 45218
rect 42364 45154 42420 45166
rect 42252 44996 42308 45006
rect 42476 44996 42532 48076
rect 42700 47124 42756 49982
rect 42812 49812 42868 49822
rect 42812 49718 42868 49756
rect 42924 49586 42980 50654
rect 44044 49924 44100 49934
rect 43260 49810 43316 49822
rect 43260 49758 43262 49810
rect 43314 49758 43316 49810
rect 43260 49700 43316 49758
rect 43260 49634 43316 49644
rect 43484 49810 43540 49822
rect 43484 49758 43486 49810
rect 43538 49758 43540 49810
rect 42924 49534 42926 49586
rect 42978 49534 42980 49586
rect 42924 49522 42980 49534
rect 43484 48356 43540 49758
rect 43932 49812 43988 49822
rect 43932 49138 43988 49756
rect 43932 49086 43934 49138
rect 43986 49086 43988 49138
rect 43932 49074 43988 49086
rect 44044 49700 44100 49868
rect 45948 49812 46004 51326
rect 46620 51266 46676 51278
rect 46620 51214 46622 51266
rect 46674 51214 46676 51266
rect 46620 50036 46676 51214
rect 48748 51266 48804 55412
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 48748 51214 48750 51266
rect 48802 51214 48804 51266
rect 48748 51202 48804 51214
rect 49532 51378 49588 51390
rect 49532 51326 49534 51378
rect 49586 51326 49588 51378
rect 48972 50370 49028 50382
rect 48972 50318 48974 50370
rect 49026 50318 49028 50370
rect 46620 49970 46676 49980
rect 47628 50036 47684 50046
rect 47628 49942 47684 49980
rect 47740 49924 47796 49934
rect 47740 49830 47796 49868
rect 45948 49746 46004 49756
rect 46956 49812 47012 49822
rect 46172 49700 46228 49710
rect 43484 48300 43764 48356
rect 42700 47058 42756 47068
rect 43036 48132 43092 48142
rect 42700 46676 42756 46686
rect 42588 46452 42644 46462
rect 42588 46358 42644 46396
rect 42252 44994 42532 44996
rect 42252 44942 42254 44994
rect 42306 44942 42532 44994
rect 42252 44940 42532 44942
rect 42252 44930 42308 44940
rect 42364 44098 42420 44110
rect 42364 44046 42366 44098
rect 42418 44046 42420 44098
rect 42364 43708 42420 44046
rect 42140 43446 42196 43484
rect 42252 43652 42420 43708
rect 42252 42980 42308 43652
rect 42140 42924 42308 42980
rect 42476 43540 42532 43550
rect 41580 42868 41636 42878
rect 41580 42774 41636 42812
rect 41580 41972 41636 41982
rect 41468 41970 41636 41972
rect 41468 41918 41582 41970
rect 41634 41918 41636 41970
rect 41468 41916 41636 41918
rect 42140 41972 42196 42924
rect 42364 42868 42420 42878
rect 42252 42756 42308 42794
rect 42364 42774 42420 42812
rect 42252 42690 42308 42700
rect 42364 41972 42420 41982
rect 42140 41970 42420 41972
rect 42140 41918 42366 41970
rect 42418 41918 42420 41970
rect 42140 41916 42420 41918
rect 41580 41906 41636 41916
rect 42364 41906 42420 41916
rect 42476 41186 42532 43484
rect 42588 42754 42644 42766
rect 42588 42702 42590 42754
rect 42642 42702 42644 42754
rect 42588 42084 42644 42702
rect 42700 42530 42756 46620
rect 43036 46562 43092 48076
rect 43708 48132 43764 48300
rect 44044 48242 44100 49644
rect 46060 49698 46228 49700
rect 46060 49646 46174 49698
rect 46226 49646 46228 49698
rect 46060 49644 46228 49646
rect 46060 49364 46116 49644
rect 46172 49634 46228 49644
rect 45836 49308 46116 49364
rect 45836 49250 45892 49308
rect 45836 49198 45838 49250
rect 45890 49198 45892 49250
rect 45836 49186 45892 49198
rect 45836 49026 45892 49038
rect 45836 48974 45838 49026
rect 45890 48974 45892 49026
rect 44716 48916 44772 48926
rect 44716 48354 44772 48860
rect 45500 48916 45556 48926
rect 45500 48822 45556 48860
rect 44716 48302 44718 48354
rect 44770 48302 44772 48354
rect 44716 48290 44772 48302
rect 44044 48190 44046 48242
rect 44098 48190 44100 48242
rect 44044 48178 44100 48190
rect 43708 48066 43764 48076
rect 44492 48132 44548 48142
rect 44492 47348 44548 48076
rect 45500 47572 45556 47582
rect 44492 47282 44548 47292
rect 45164 47570 45556 47572
rect 45164 47518 45502 47570
rect 45554 47518 45556 47570
rect 45164 47516 45556 47518
rect 45164 46786 45220 47516
rect 45500 47506 45556 47516
rect 45612 47348 45668 47358
rect 45612 47254 45668 47292
rect 45836 47346 45892 48974
rect 46956 48804 47012 49756
rect 48972 49812 49028 50318
rect 48972 49746 49028 49756
rect 49532 49812 49588 51326
rect 50316 51266 50372 51278
rect 50316 51214 50318 51266
rect 50370 51214 50372 51266
rect 50316 50482 50372 51214
rect 52444 51268 52500 51278
rect 52444 51174 52500 51212
rect 53004 51266 53060 51278
rect 53004 51214 53006 51266
rect 53058 51214 53060 51266
rect 50316 50430 50318 50482
rect 50370 50430 50372 50482
rect 50316 50418 50372 50430
rect 53004 50372 53060 51214
rect 55132 51268 55188 51278
rect 53340 50484 53396 50494
rect 53340 50372 53396 50428
rect 54236 50484 54292 50494
rect 54236 50390 54292 50428
rect 53004 50370 53396 50372
rect 53004 50318 53342 50370
rect 53394 50318 53396 50370
rect 53004 50316 53396 50318
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 47516 49586 47572 49598
rect 47516 49534 47518 49586
rect 47570 49534 47572 49586
rect 47180 48804 47236 48814
rect 46956 48802 47236 48804
rect 46956 48750 47182 48802
rect 47234 48750 47236 48802
rect 46956 48748 47236 48750
rect 47180 47460 47236 48748
rect 45836 47294 45838 47346
rect 45890 47294 45892 47346
rect 45836 47236 45892 47294
rect 45836 47170 45892 47180
rect 46956 47458 47236 47460
rect 46956 47406 47182 47458
rect 47234 47406 47236 47458
rect 46956 47404 47236 47406
rect 45164 46734 45166 46786
rect 45218 46734 45220 46786
rect 45164 46722 45220 46734
rect 43036 46510 43038 46562
rect 43090 46510 43092 46562
rect 43036 46498 43092 46510
rect 45836 46676 45892 46686
rect 46396 46676 46452 46686
rect 46956 46676 47012 47404
rect 47180 47394 47236 47404
rect 47180 47236 47236 47246
rect 47180 46898 47236 47180
rect 47516 47236 47572 49534
rect 49532 49026 49588 49756
rect 51100 49812 51156 49822
rect 51100 49718 51156 49756
rect 53004 49812 53060 50316
rect 53340 50306 53396 50316
rect 53004 49746 53060 49756
rect 53564 49812 53620 49822
rect 51884 49700 51940 49710
rect 51884 49698 52052 49700
rect 51884 49646 51886 49698
rect 51938 49646 52052 49698
rect 51884 49644 52052 49646
rect 51884 49634 51940 49644
rect 49532 48974 49534 49026
rect 49586 48974 49588 49026
rect 49532 48962 49588 48974
rect 48972 48916 49028 48926
rect 48972 48822 49028 48860
rect 50316 48916 50372 48926
rect 50316 48822 50372 48860
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 48076 48354 48132 48366
rect 48076 48302 48078 48354
rect 48130 48302 48132 48354
rect 47964 47572 48020 47582
rect 48076 47572 48132 48302
rect 48748 48244 48804 48254
rect 48748 48150 48804 48188
rect 49532 48244 49588 48254
rect 49532 48150 49588 48188
rect 50876 48244 50932 48254
rect 47964 47570 48132 47572
rect 47964 47518 47966 47570
rect 48018 47518 48132 47570
rect 47964 47516 48132 47518
rect 50092 47572 50148 47582
rect 47964 47506 48020 47516
rect 50092 47478 50148 47516
rect 50540 47236 50596 47246
rect 47516 47170 47572 47180
rect 50428 47234 50596 47236
rect 50428 47182 50542 47234
rect 50594 47182 50596 47234
rect 50428 47180 50596 47182
rect 47180 46846 47182 46898
rect 47234 46846 47236 46898
rect 47180 46834 47236 46846
rect 48412 46788 48468 46798
rect 45836 46674 47012 46676
rect 45836 46622 45838 46674
rect 45890 46622 46398 46674
rect 46450 46622 47012 46674
rect 45836 46620 47012 46622
rect 43932 46002 43988 46014
rect 43932 45950 43934 46002
rect 43986 45950 43988 46002
rect 43820 45892 43876 45902
rect 43820 45108 43876 45836
rect 43932 45444 43988 45950
rect 45612 45892 45668 45902
rect 45836 45892 45892 46620
rect 46396 46610 46452 46620
rect 46956 46004 47012 46620
rect 47068 46674 47124 46686
rect 47068 46622 47070 46674
rect 47122 46622 47124 46674
rect 47068 46452 47124 46622
rect 47740 46674 47796 46686
rect 47740 46622 47742 46674
rect 47794 46622 47796 46674
rect 47740 46564 47796 46622
rect 48412 46674 48468 46732
rect 48412 46622 48414 46674
rect 48466 46622 48468 46674
rect 48412 46610 48468 46622
rect 48524 46786 48580 46798
rect 48524 46734 48526 46786
rect 48578 46734 48580 46786
rect 47740 46498 47796 46508
rect 47068 46386 47124 46396
rect 46956 45938 47012 45948
rect 48412 46002 48468 46014
rect 48412 45950 48414 46002
rect 48466 45950 48468 46002
rect 45612 45890 45892 45892
rect 45612 45838 45614 45890
rect 45666 45838 45892 45890
rect 45612 45836 45892 45838
rect 45612 45826 45668 45836
rect 46284 45778 46340 45790
rect 46284 45726 46286 45778
rect 46338 45726 46340 45778
rect 43932 45378 43988 45388
rect 44380 45666 44436 45678
rect 44380 45614 44382 45666
rect 44434 45614 44436 45666
rect 44380 45108 44436 45614
rect 43820 45106 44436 45108
rect 43820 45054 43822 45106
rect 43874 45054 44436 45106
rect 43820 45052 44436 45054
rect 42812 42754 42868 42766
rect 42812 42702 42814 42754
rect 42866 42702 42868 42754
rect 42812 42644 42868 42702
rect 43820 42756 43876 45052
rect 44492 44994 44548 45006
rect 44492 44942 44494 44994
rect 44546 44942 44548 44994
rect 44492 44212 44548 44942
rect 44604 44212 44660 44222
rect 44492 44210 44660 44212
rect 44492 44158 44606 44210
rect 44658 44158 44660 44210
rect 44492 44156 44660 44158
rect 46284 44212 46340 45726
rect 46620 44996 46676 45006
rect 46620 44902 46676 44940
rect 47068 44994 47124 45006
rect 47068 44942 47070 44994
rect 47122 44942 47124 44994
rect 46396 44212 46452 44222
rect 46284 44210 46452 44212
rect 46284 44158 46398 44210
rect 46450 44158 46452 44210
rect 46284 44156 46452 44158
rect 44604 44146 44660 44156
rect 46396 44146 46452 44156
rect 45836 44098 45892 44110
rect 45836 44046 45838 44098
rect 45890 44046 45892 44098
rect 45836 43708 45892 44046
rect 45836 43652 46340 43708
rect 46284 42866 46340 43652
rect 46284 42814 46286 42866
rect 46338 42814 46340 42866
rect 46284 42802 46340 42814
rect 46956 43652 47012 43662
rect 47068 43652 47124 44942
rect 47404 44996 47460 45006
rect 47404 44210 47460 44940
rect 47404 44158 47406 44210
rect 47458 44158 47460 44210
rect 47404 44146 47460 44158
rect 48076 44322 48132 44334
rect 48076 44270 48078 44322
rect 48130 44270 48132 44322
rect 48076 43708 48132 44270
rect 48412 44212 48468 45950
rect 48524 44434 48580 46734
rect 50428 46676 50484 47180
rect 50540 47170 50596 47180
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 49532 46564 49588 46574
rect 49532 46470 49588 46508
rect 48972 46004 49028 46014
rect 48972 45910 49028 45948
rect 50428 46004 50484 46620
rect 50428 45938 50484 45948
rect 49756 45668 49812 45678
rect 49756 45666 50372 45668
rect 49756 45614 49758 45666
rect 49810 45614 50372 45666
rect 49756 45612 50372 45614
rect 49756 45602 49812 45612
rect 50316 45218 50372 45612
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50316 45166 50318 45218
rect 50370 45166 50372 45218
rect 50316 45154 50372 45166
rect 48524 44382 48526 44434
rect 48578 44382 48580 44434
rect 48524 44370 48580 44382
rect 49644 45106 49700 45118
rect 49644 45054 49646 45106
rect 49698 45054 49700 45106
rect 49084 44322 49140 44334
rect 49084 44270 49086 44322
rect 49138 44270 49140 44322
rect 48412 44146 48468 44156
rect 48972 44212 49028 44222
rect 48972 44118 49028 44156
rect 48412 43764 48468 43802
rect 49084 43708 49140 44270
rect 48076 43652 48356 43708
rect 48412 43698 48468 43708
rect 46956 43650 47124 43652
rect 46956 43598 46958 43650
rect 47010 43598 47124 43650
rect 46956 43596 47124 43598
rect 43820 42690 43876 42700
rect 44716 42756 44772 42766
rect 44716 42662 44772 42700
rect 44940 42756 44996 42766
rect 42812 42578 42868 42588
rect 44492 42644 44548 42654
rect 42700 42478 42702 42530
rect 42754 42478 42756 42530
rect 42700 42466 42756 42478
rect 42588 42018 42644 42028
rect 44492 41858 44548 42588
rect 44940 42194 44996 42700
rect 45612 42756 45668 42766
rect 45612 42662 45668 42700
rect 46956 42756 47012 43596
rect 48300 42868 48356 43652
rect 48972 43652 49140 43708
rect 48412 42868 48468 42878
rect 48300 42866 48468 42868
rect 48300 42814 48414 42866
rect 48466 42814 48468 42866
rect 48300 42812 48468 42814
rect 48412 42802 48468 42812
rect 48972 42866 49028 43652
rect 49420 43428 49476 43438
rect 49420 43334 49476 43372
rect 48972 42814 48974 42866
rect 49026 42814 49028 42866
rect 48972 42802 49028 42814
rect 46956 42690 47012 42700
rect 44940 42142 44942 42194
rect 44994 42142 44996 42194
rect 44940 42130 44996 42142
rect 49644 42084 49700 45054
rect 50876 44434 50932 48188
rect 51548 48130 51604 48142
rect 51548 48078 51550 48130
rect 51602 48078 51604 48130
rect 51548 47012 51604 48078
rect 51996 47348 52052 49644
rect 52444 49138 52500 49150
rect 52444 49086 52446 49138
rect 52498 49086 52500 49138
rect 52444 47460 52500 49086
rect 53564 49026 53620 49756
rect 54012 49698 54068 49710
rect 54012 49646 54014 49698
rect 54066 49646 54068 49698
rect 54012 49140 54068 49646
rect 54012 49084 54628 49140
rect 53564 48974 53566 49026
rect 53618 48974 53620 49026
rect 53564 48962 53620 48974
rect 54348 48916 54404 48926
rect 52444 47394 52500 47404
rect 53452 47572 53508 47582
rect 52108 47348 52164 47358
rect 51996 47346 52164 47348
rect 51996 47294 52110 47346
rect 52162 47294 52164 47346
rect 51996 47292 52164 47294
rect 52108 47282 52164 47292
rect 53452 47346 53508 47516
rect 54012 47460 54068 47470
rect 54012 47366 54068 47404
rect 53452 47294 53454 47346
rect 53506 47294 53508 47346
rect 53452 47282 53508 47294
rect 52668 47234 52724 47246
rect 52668 47182 52670 47234
rect 52722 47182 52724 47234
rect 52668 47124 52724 47182
rect 52668 47058 52724 47068
rect 54012 47234 54068 47246
rect 54012 47182 54014 47234
rect 54066 47182 54068 47234
rect 51212 46676 51268 46686
rect 51212 46582 51268 46620
rect 51548 46676 51604 46956
rect 54012 46788 54068 47182
rect 54012 46722 54068 46732
rect 54348 46676 54404 48860
rect 54572 47348 54628 49084
rect 55132 47458 55188 51212
rect 56140 49812 56196 49822
rect 56140 49810 56532 49812
rect 56140 49758 56142 49810
rect 56194 49758 56532 49810
rect 56140 49756 56532 49758
rect 56140 49746 56196 49756
rect 55356 49698 55412 49710
rect 55356 49646 55358 49698
rect 55410 49646 55412 49698
rect 55356 49140 55412 49646
rect 55356 49074 55412 49084
rect 56476 49138 56532 49756
rect 56476 49086 56478 49138
rect 56530 49086 56532 49138
rect 56476 49074 56532 49086
rect 56924 48916 56980 48926
rect 56924 48822 56980 48860
rect 55132 47406 55134 47458
rect 55186 47406 55188 47458
rect 55132 47394 55188 47406
rect 55020 47348 55076 47358
rect 54572 47346 55076 47348
rect 54572 47294 55022 47346
rect 55074 47294 55076 47346
rect 54572 47292 55076 47294
rect 55020 47282 55076 47292
rect 54572 47012 54628 47022
rect 54572 46898 54628 46956
rect 54572 46846 54574 46898
rect 54626 46846 54628 46898
rect 54572 46834 54628 46846
rect 54348 46620 54628 46676
rect 51548 46610 51604 46620
rect 51996 46562 52052 46574
rect 51996 46510 51998 46562
rect 52050 46510 52052 46562
rect 51996 45780 52052 46510
rect 54124 46562 54180 46574
rect 54124 46510 54126 46562
rect 54178 46510 54180 46562
rect 52108 45780 52164 45790
rect 51996 45778 52164 45780
rect 51996 45726 52110 45778
rect 52162 45726 52164 45778
rect 51996 45724 52164 45726
rect 52108 45714 52164 45724
rect 54012 45668 54068 45678
rect 53788 45666 54068 45668
rect 53788 45614 54014 45666
rect 54066 45614 54068 45666
rect 53788 45612 54068 45614
rect 53788 45218 53844 45612
rect 54012 45602 54068 45612
rect 53788 45166 53790 45218
rect 53842 45166 53844 45218
rect 53788 45154 53844 45166
rect 53004 45108 53060 45118
rect 52668 45106 53060 45108
rect 52668 45054 53006 45106
rect 53058 45054 53060 45106
rect 52668 45052 53060 45054
rect 50876 44382 50878 44434
rect 50930 44382 50932 44434
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50652 43652 50708 43662
rect 50428 43650 50708 43652
rect 50428 43598 50654 43650
rect 50706 43598 50708 43650
rect 50428 43596 50708 43598
rect 50428 42196 50484 43596
rect 50652 43586 50708 43596
rect 50876 43428 50932 44382
rect 52444 44994 52500 45006
rect 52444 44942 52446 44994
rect 52498 44942 52500 44994
rect 52444 44324 52500 44942
rect 52668 44434 52724 45052
rect 52668 44382 52670 44434
rect 52722 44382 52724 44434
rect 52668 44370 52724 44382
rect 52444 44258 52500 44268
rect 50876 43362 50932 43372
rect 51100 43764 51156 43774
rect 51100 42866 51156 43708
rect 52332 43652 52388 43662
rect 51100 42814 51102 42866
rect 51154 42814 51156 42866
rect 51100 42802 51156 42814
rect 51212 43538 51268 43550
rect 51212 43486 51214 43538
rect 51266 43486 51268 43538
rect 51212 43428 51268 43486
rect 50876 42756 50932 42766
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50428 42140 50820 42196
rect 49644 42018 49700 42028
rect 50092 42084 50148 42094
rect 50092 41970 50148 42028
rect 50092 41918 50094 41970
rect 50146 41918 50148 41970
rect 50092 41906 50148 41918
rect 50764 41970 50820 42140
rect 50764 41918 50766 41970
rect 50818 41918 50820 41970
rect 50764 41906 50820 41918
rect 50876 42084 50932 42700
rect 44492 41806 44494 41858
rect 44546 41806 44548 41858
rect 44492 41794 44548 41806
rect 42476 41134 42478 41186
rect 42530 41134 42532 41186
rect 40684 40238 40686 40290
rect 40738 40238 40740 40290
rect 40684 40226 40740 40238
rect 40908 41074 40964 41086
rect 40908 41022 40910 41074
rect 40962 41022 40964 41074
rect 40908 40404 40964 41022
rect 42476 40964 42532 41134
rect 42476 40898 42532 40908
rect 44380 40964 44436 40974
rect 44380 40870 44436 40908
rect 46844 40964 46900 40974
rect 40908 39618 40964 40348
rect 46620 40402 46676 40414
rect 46620 40350 46622 40402
rect 46674 40350 46676 40402
rect 43708 40292 43764 40302
rect 45836 40292 45892 40302
rect 43708 40290 44660 40292
rect 43708 40238 43710 40290
rect 43762 40238 44660 40290
rect 43708 40236 44660 40238
rect 43708 40226 43764 40236
rect 43820 39732 43876 39742
rect 43820 39730 44212 39732
rect 43820 39678 43822 39730
rect 43874 39678 44212 39730
rect 43820 39676 44212 39678
rect 43820 39666 43876 39676
rect 40908 39566 40910 39618
rect 40962 39566 40964 39618
rect 40908 39554 40964 39566
rect 41692 39508 41748 39518
rect 41692 39506 41972 39508
rect 41692 39454 41694 39506
rect 41746 39454 41972 39506
rect 41692 39452 41972 39454
rect 41692 39442 41748 39452
rect 40012 39342 40014 39394
rect 40066 39342 40068 39394
rect 40012 38836 40068 39342
rect 41916 39058 41972 39452
rect 41916 39006 41918 39058
rect 41970 39006 41972 39058
rect 41916 38994 41972 39006
rect 43372 39060 43428 39070
rect 43372 38966 43428 39004
rect 44044 39060 44100 39070
rect 44044 38966 44100 39004
rect 40572 38948 40628 38958
rect 40572 38946 41860 38948
rect 40572 38894 40574 38946
rect 40626 38894 41860 38946
rect 40572 38892 41860 38894
rect 40572 38882 40628 38892
rect 40012 38770 40068 38780
rect 40348 38724 40404 38734
rect 37660 38546 37716 38556
rect 39676 38612 39732 38622
rect 37548 38164 37604 38174
rect 37548 38070 37604 38108
rect 39676 38162 39732 38556
rect 39676 38110 39678 38162
rect 39730 38110 39732 38162
rect 39676 38098 39732 38110
rect 40348 38052 40404 38668
rect 41804 38162 41860 38892
rect 42924 38834 42980 38846
rect 43148 38836 43204 38846
rect 42924 38782 42926 38834
rect 42978 38782 42980 38834
rect 41804 38110 41806 38162
rect 41858 38110 41860 38162
rect 41804 38098 41860 38110
rect 42812 38724 42868 38734
rect 41020 38052 41076 38062
rect 40348 38050 41524 38052
rect 40348 37998 40350 38050
rect 40402 37998 41022 38050
rect 41074 37998 41524 38050
rect 40348 37996 41524 37998
rect 40348 37986 40404 37996
rect 37884 37940 37940 37950
rect 37324 37214 37326 37266
rect 37378 37214 37380 37266
rect 37324 37202 37380 37214
rect 37436 37378 37492 37390
rect 37436 37326 37438 37378
rect 37490 37326 37492 37378
rect 37436 37156 37492 37326
rect 37436 37090 37492 37100
rect 37660 37266 37716 37278
rect 37660 37214 37662 37266
rect 37714 37214 37716 37266
rect 36988 36530 37044 36540
rect 37548 36596 37604 36606
rect 37548 36502 37604 36540
rect 33068 35588 33124 35598
rect 33068 34916 33124 35532
rect 36092 35588 36148 35598
rect 36092 35494 36148 35532
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 32172 34018 32340 34020
rect 32172 33966 32174 34018
rect 32226 33966 32340 34018
rect 32172 33964 32340 33966
rect 32620 34914 33124 34916
rect 32620 34862 33070 34914
rect 33122 34862 33124 34914
rect 32620 34860 33124 34862
rect 32620 34354 32676 34860
rect 33068 34850 33124 34860
rect 35868 35026 35924 35038
rect 35868 34974 35870 35026
rect 35922 34974 35924 35026
rect 32620 34302 32622 34354
rect 32674 34302 32676 34354
rect 32172 33954 32228 33964
rect 32620 33458 32676 34302
rect 33740 34802 33796 34814
rect 33740 34750 33742 34802
rect 33794 34750 33796 34802
rect 33740 34356 33796 34750
rect 33852 34356 33908 34366
rect 33740 34354 33908 34356
rect 33740 34302 33854 34354
rect 33906 34302 33908 34354
rect 33740 34300 33908 34302
rect 33852 34290 33908 34300
rect 35308 34020 35364 34030
rect 35308 33926 35364 33964
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 32620 33406 32622 33458
rect 32674 33406 32676 33458
rect 29596 32788 29652 32798
rect 28364 32622 28366 32674
rect 28418 32622 28420 32674
rect 28364 32610 28420 32622
rect 29148 32786 29764 32788
rect 29148 32734 29598 32786
rect 29650 32734 29764 32786
rect 29148 32732 29764 32734
rect 29148 32562 29204 32732
rect 29596 32722 29652 32732
rect 29148 32510 29150 32562
rect 29202 32510 29204 32562
rect 29148 32498 29204 32510
rect 27020 32452 27076 32462
rect 26572 31892 26852 31948
rect 26348 30996 26404 31006
rect 26236 30994 26404 30996
rect 26236 30942 26350 30994
rect 26402 30942 26404 30994
rect 26236 30940 26404 30942
rect 26348 30930 26404 30940
rect 26796 30994 26852 31892
rect 26796 30942 26798 30994
rect 26850 30942 26852 30994
rect 26796 30930 26852 30942
rect 26908 31890 26964 31902
rect 26908 31838 26910 31890
rect 26962 31838 26964 31890
rect 24780 30046 24782 30098
rect 24834 30046 24836 30098
rect 24780 30034 24836 30046
rect 26236 30770 26292 30782
rect 26236 30718 26238 30770
rect 26290 30718 26292 30770
rect 24108 29362 24164 29372
rect 24892 29314 24948 29326
rect 24892 29262 24894 29314
rect 24946 29262 24948 29314
rect 24892 28868 24948 29262
rect 24892 28802 24948 28812
rect 25900 28868 25956 28878
rect 25900 28774 25956 28812
rect 21756 28702 21758 28754
rect 21810 28702 21812 28754
rect 21756 28690 21812 28702
rect 25676 28642 25732 28654
rect 25676 28590 25678 28642
rect 25730 28590 25732 28642
rect 21196 28420 21252 28430
rect 20748 27806 20750 27858
rect 20802 27806 20804 27858
rect 20748 27794 20804 27806
rect 20860 27970 20916 27982
rect 20860 27918 20862 27970
rect 20914 27918 20916 27970
rect 15820 27746 15876 27758
rect 15820 27694 15822 27746
rect 15874 27694 15876 27746
rect 15820 27300 15876 27694
rect 16380 27748 16436 27758
rect 16380 27654 16436 27692
rect 15820 27234 15876 27244
rect 18284 26852 18340 26862
rect 18284 26850 18564 26852
rect 18284 26798 18286 26850
rect 18338 26798 18564 26850
rect 18284 26796 18564 26798
rect 18284 26786 18340 26796
rect 18508 26402 18564 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 18508 26350 18510 26402
rect 18562 26350 18564 26402
rect 18508 26338 18564 26350
rect 17836 26290 17892 26302
rect 17836 26238 17838 26290
rect 17890 26238 17892 26290
rect 15820 25508 15876 25518
rect 15820 25414 15876 25452
rect 17836 25508 17892 26238
rect 20636 26178 20692 26190
rect 20636 26126 20638 26178
rect 20690 26126 20692 26178
rect 20524 25732 20580 25742
rect 20636 25732 20692 26126
rect 20524 25730 20692 25732
rect 20524 25678 20526 25730
rect 20578 25678 20692 25730
rect 20524 25676 20692 25678
rect 20860 25730 20916 27918
rect 21196 27970 21252 28364
rect 25116 28420 25172 28430
rect 25116 28418 25620 28420
rect 25116 28366 25118 28418
rect 25170 28366 25620 28418
rect 25116 28364 25620 28366
rect 25116 28354 25172 28364
rect 21756 28084 21812 28094
rect 21756 27990 21812 28028
rect 21196 27918 21198 27970
rect 21250 27918 21252 27970
rect 21196 27906 21252 27918
rect 21532 27972 21588 27982
rect 22540 27972 22596 27982
rect 21532 27858 21588 27916
rect 21532 27806 21534 27858
rect 21586 27806 21588 27858
rect 21532 27794 21588 27806
rect 22316 27970 22596 27972
rect 22316 27918 22542 27970
rect 22594 27918 22596 27970
rect 22316 27916 22596 27918
rect 20860 25678 20862 25730
rect 20914 25678 20916 25730
rect 20524 25666 20580 25676
rect 20860 25666 20916 25678
rect 20972 26962 21028 26974
rect 20972 26910 20974 26962
rect 21026 26910 21028 26962
rect 18620 25620 18676 25630
rect 18620 25526 18676 25564
rect 20300 25620 20356 25630
rect 17836 25442 17892 25452
rect 18284 25508 18340 25518
rect 16492 25394 16548 25406
rect 16492 25342 16494 25394
rect 16546 25342 16548 25394
rect 16492 24948 16548 25342
rect 16492 24882 16548 24892
rect 17724 24948 17780 24958
rect 17724 24854 17780 24892
rect 18284 24610 18340 25452
rect 20188 25508 20244 25546
rect 20300 25526 20356 25564
rect 20188 25442 20244 25452
rect 20748 25506 20804 25518
rect 20748 25454 20750 25506
rect 20802 25454 20804 25506
rect 19516 25282 19572 25294
rect 19516 25230 19518 25282
rect 19570 25230 19572 25282
rect 19516 24836 19572 25230
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19628 24836 19684 24846
rect 19516 24834 19684 24836
rect 19516 24782 19630 24834
rect 19682 24782 19684 24834
rect 19516 24780 19684 24782
rect 19628 24770 19684 24780
rect 18284 24558 18286 24610
rect 18338 24558 18340 24610
rect 16604 24050 16660 24062
rect 16604 23998 16606 24050
rect 16658 23998 16660 24050
rect 16604 23604 16660 23998
rect 17052 24052 17108 24062
rect 17052 23958 17108 23996
rect 16604 23538 16660 23548
rect 17948 23716 18004 23726
rect 16604 23380 16660 23390
rect 16604 23286 16660 23324
rect 15372 23212 15652 23268
rect 15260 23100 15540 23156
rect 15484 23042 15540 23100
rect 15484 22990 15486 23042
rect 15538 22990 15540 23042
rect 15484 22978 15540 22990
rect 15260 22484 15316 22494
rect 15260 22390 15316 22428
rect 13132 21758 13134 21810
rect 13186 21758 13188 21810
rect 13132 21588 13188 21758
rect 14140 22370 14644 22372
rect 14140 22318 14590 22370
rect 14642 22318 14644 22370
rect 14140 22316 14644 22318
rect 14140 21810 14196 22316
rect 14588 22306 14644 22316
rect 14140 21758 14142 21810
rect 14194 21758 14196 21810
rect 14140 21746 14196 21758
rect 13132 21522 13188 21532
rect 13468 20580 13524 20590
rect 12796 20132 13300 20188
rect 12572 19348 12628 19358
rect 12572 19254 12628 19292
rect 13244 18562 13300 20132
rect 13468 19348 13524 20524
rect 14812 20578 14868 20590
rect 14812 20526 14814 20578
rect 14866 20526 14868 20578
rect 14700 20132 14756 20142
rect 14812 20132 14868 20526
rect 14700 20130 14868 20132
rect 14700 20078 14702 20130
rect 14754 20078 14868 20130
rect 14700 20076 14868 20078
rect 15484 20578 15540 20590
rect 15484 20526 15486 20578
rect 15538 20526 15540 20578
rect 14700 20066 14756 20076
rect 14028 20018 14084 20030
rect 14028 19966 14030 20018
rect 14082 19966 14084 20018
rect 13580 19348 13636 19358
rect 13244 18510 13246 18562
rect 13298 18510 13300 18562
rect 13244 18498 13300 18510
rect 13356 19346 13636 19348
rect 13356 19294 13582 19346
rect 13634 19294 13636 19346
rect 13356 19292 13636 19294
rect 13132 18450 13188 18462
rect 13132 18398 13134 18450
rect 13186 18398 13188 18450
rect 12684 18228 12740 18238
rect 11788 17714 11844 17724
rect 12572 18226 12740 18228
rect 12572 18174 12686 18226
rect 12738 18174 12740 18226
rect 12572 18172 12740 18174
rect 9660 16818 9716 16828
rect 9772 16994 9828 17006
rect 9772 16942 9774 16994
rect 9826 16942 9828 16994
rect 8764 16098 8820 16716
rect 9436 16212 9492 16222
rect 9772 16212 9828 16942
rect 10780 16884 10836 16894
rect 10780 16790 10836 16828
rect 11452 16884 11508 16894
rect 11452 16790 11508 16828
rect 12124 16770 12180 16782
rect 12124 16718 12126 16770
rect 12178 16718 12180 16770
rect 9436 16210 9828 16212
rect 9436 16158 9438 16210
rect 9490 16158 9828 16210
rect 9436 16156 9828 16158
rect 11564 16212 11620 16222
rect 9436 16146 9492 16156
rect 11564 16118 11620 16156
rect 8764 16046 8766 16098
rect 8818 16046 8820 16098
rect 8764 15092 8820 16046
rect 12124 15988 12180 16718
rect 12236 15988 12292 15998
rect 12124 15986 12292 15988
rect 12124 15934 12238 15986
rect 12290 15934 12292 15986
rect 12124 15932 12292 15934
rect 12236 15922 12292 15932
rect 10108 15204 10164 15214
rect 10108 15202 10836 15204
rect 10108 15150 10110 15202
rect 10162 15150 10836 15202
rect 10108 15148 10836 15150
rect 10108 15138 10164 15148
rect 8764 15026 8820 15036
rect 9996 15090 10052 15102
rect 9996 15038 9998 15090
rect 10050 15038 10052 15090
rect 8652 14420 8708 14430
rect 8652 14418 9268 14420
rect 8652 14366 8654 14418
rect 8706 14366 9268 14418
rect 8652 14364 9268 14366
rect 8652 14354 8708 14364
rect 8652 13860 8708 13870
rect 8428 13858 8708 13860
rect 8428 13806 8654 13858
rect 8706 13806 8708 13858
rect 8428 13804 8708 13806
rect 8652 13748 8708 13804
rect 8652 13682 8708 13692
rect 8988 13860 9044 13870
rect 8988 13746 9044 13804
rect 8988 13694 8990 13746
rect 9042 13694 9044 13746
rect 8988 13682 9044 13694
rect 8988 12964 9044 12974
rect 8988 12870 9044 12908
rect 9100 12852 9156 12862
rect 9100 12758 9156 12796
rect 9212 12738 9268 14364
rect 9996 13972 10052 15038
rect 10780 14642 10836 15148
rect 10780 14590 10782 14642
rect 10834 14590 10836 14642
rect 10780 14578 10836 14590
rect 11340 15092 11396 15102
rect 11340 14642 11396 15036
rect 11340 14590 11342 14642
rect 11394 14590 11396 14642
rect 11340 14578 11396 14590
rect 9996 13916 10948 13972
rect 9996 13748 10052 13758
rect 9996 13654 10052 13692
rect 10220 13634 10276 13646
rect 10220 13582 10222 13634
rect 10274 13582 10276 13634
rect 9212 12686 9214 12738
rect 9266 12686 9268 12738
rect 9212 12674 9268 12686
rect 9548 12962 9604 12974
rect 9548 12910 9550 12962
rect 9602 12910 9604 12962
rect 8316 12114 8372 12124
rect 8988 12180 9044 12190
rect 8204 11330 8260 11340
rect 8652 11506 8708 11518
rect 8652 11454 8654 11506
rect 8706 11454 8708 11506
rect 6972 10610 7308 10612
rect 6972 10558 6974 10610
rect 7026 10558 7308 10610
rect 6972 10556 7308 10558
rect 6972 10546 7028 10556
rect 3948 10500 4004 10510
rect 7308 10480 7364 10556
rect 7420 10610 7476 10622
rect 7420 10558 7422 10610
rect 7474 10558 7476 10610
rect 3948 10406 4004 10444
rect 2604 9886 2606 9938
rect 2658 9886 2660 9938
rect 2604 9874 2660 9886
rect 3052 9884 3220 9940
rect 3276 10332 3444 10388
rect 7196 10386 7252 10398
rect 7196 10334 7198 10386
rect 7250 10334 7252 10386
rect 3052 8428 3108 9884
rect 3276 8930 3332 10332
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4732 9938 4788 9950
rect 4732 9886 4734 9938
rect 4786 9886 4788 9938
rect 4732 9716 4788 9886
rect 7196 9940 7252 10334
rect 7196 9874 7252 9884
rect 6972 9828 7028 9838
rect 6972 9734 7028 9772
rect 3276 8878 3278 8930
rect 3330 8878 3332 8930
rect 3276 8866 3332 8878
rect 3388 9156 3444 9166
rect 3388 8930 3444 9100
rect 4060 9044 4116 9054
rect 4060 8950 4116 8988
rect 4732 9044 4788 9660
rect 6748 9716 6804 9726
rect 6748 9622 6804 9660
rect 6860 9714 6916 9726
rect 6860 9662 6862 9714
rect 6914 9662 6916 9714
rect 6860 9492 6916 9662
rect 5964 9156 6020 9166
rect 5964 9062 6020 9100
rect 6860 9156 6916 9436
rect 6860 9090 6916 9100
rect 7196 9716 7252 9726
rect 4732 8978 4788 8988
rect 4956 9044 5012 9054
rect 3388 8878 3390 8930
rect 3442 8878 3444 8930
rect 3388 8428 3444 8878
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 2940 8372 3108 8428
rect 3164 8372 3444 8428
rect 2828 8146 2884 8158
rect 2828 8094 2830 8146
rect 2882 8094 2884 8146
rect 2828 7698 2884 8094
rect 2828 7646 2830 7698
rect 2882 7646 2884 7698
rect 2828 7634 2884 7646
rect 2604 7476 2660 7486
rect 2828 7476 2884 7486
rect 2940 7476 2996 8372
rect 3164 7586 3220 8372
rect 4956 8370 5012 8988
rect 6188 9044 6244 9054
rect 6188 8950 6244 8988
rect 7196 9042 7252 9660
rect 7420 9604 7476 10558
rect 8204 10612 8260 10622
rect 8092 9940 8148 9950
rect 8092 9846 8148 9884
rect 7420 9510 7476 9548
rect 7868 9826 7924 9838
rect 7868 9774 7870 9826
rect 7922 9774 7924 9826
rect 7868 9492 7924 9774
rect 7868 9426 7924 9436
rect 8204 9266 8260 10556
rect 8540 9828 8596 9838
rect 8652 9828 8708 11454
rect 8988 11172 9044 12124
rect 9548 11956 9604 12910
rect 9772 12404 9828 12414
rect 9772 12310 9828 12348
rect 9548 11890 9604 11900
rect 10108 11956 10164 11966
rect 10108 11862 10164 11900
rect 10220 11620 10276 13582
rect 10332 12852 10388 13916
rect 10444 13748 10500 13758
rect 10444 13654 10500 13692
rect 10892 13746 10948 13916
rect 10892 13694 10894 13746
rect 10946 13694 10948 13746
rect 10892 13682 10948 13694
rect 12572 13748 12628 18172
rect 12684 18162 12740 18172
rect 13132 18228 13188 18398
rect 13132 18162 13188 18172
rect 13356 17892 13412 19292
rect 13580 19282 13636 19292
rect 13916 19348 13972 19358
rect 12684 17836 13412 17892
rect 13468 18450 13524 18462
rect 13468 18398 13470 18450
rect 13522 18398 13524 18450
rect 12684 17778 12740 17836
rect 12684 17726 12686 17778
rect 12738 17726 12740 17778
rect 12684 17714 12740 17726
rect 12796 16772 12852 17836
rect 12796 16210 12852 16716
rect 12796 16158 12798 16210
rect 12850 16158 12852 16210
rect 12796 16146 12852 16158
rect 13468 15876 13524 18398
rect 13580 17780 13636 17790
rect 13580 17686 13636 17724
rect 13916 16322 13972 19292
rect 14028 18452 14084 19966
rect 14140 18452 14196 18462
rect 14028 18396 14140 18452
rect 14140 18358 14196 18396
rect 14812 18340 14868 18350
rect 14812 18246 14868 18284
rect 15484 18340 15540 20526
rect 15596 19348 15652 23212
rect 16044 23266 16100 23278
rect 16044 23214 16046 23266
rect 16098 23214 16100 23266
rect 16044 22484 16100 23214
rect 16044 22418 16100 22428
rect 17388 22484 17444 22494
rect 17388 22390 17444 22428
rect 17948 22370 18004 23660
rect 18284 23716 18340 24558
rect 18284 23650 18340 23660
rect 18844 24722 18900 24734
rect 18844 24670 18846 24722
rect 18898 24670 18900 24722
rect 18844 23716 18900 24670
rect 20748 24612 20804 25454
rect 20748 24546 20804 24556
rect 20860 25508 20916 25518
rect 18844 23650 18900 23660
rect 18956 23714 19012 23726
rect 18956 23662 18958 23714
rect 19010 23662 19012 23714
rect 18508 23604 18564 23614
rect 17948 22318 17950 22370
rect 18002 22318 18004 22370
rect 17948 20802 18004 22318
rect 17948 20750 17950 20802
rect 18002 20750 18004 20802
rect 17052 20580 17108 20590
rect 17948 20580 18004 20750
rect 17052 20578 18004 20580
rect 17052 20526 17054 20578
rect 17106 20526 18004 20578
rect 17052 20524 18004 20526
rect 18060 22484 18116 22494
rect 16828 19908 16884 19918
rect 16828 19814 16884 19852
rect 15596 19234 15652 19292
rect 15596 19182 15598 19234
rect 15650 19182 15652 19234
rect 15596 19170 15652 19182
rect 16940 19796 16996 19806
rect 15484 18274 15540 18284
rect 16604 18452 16660 18462
rect 14924 16996 14980 17006
rect 14924 16994 15092 16996
rect 14924 16942 14926 16994
rect 14978 16942 15092 16994
rect 14924 16940 15092 16942
rect 14924 16930 14980 16940
rect 14252 16770 14308 16782
rect 14252 16718 14254 16770
rect 14306 16718 14308 16770
rect 13916 16270 13918 16322
rect 13970 16270 13972 16322
rect 13916 16258 13972 16270
rect 14140 16324 14196 16334
rect 14252 16324 14308 16718
rect 14140 16322 14308 16324
rect 14140 16270 14142 16322
rect 14194 16270 14308 16322
rect 14140 16268 14308 16270
rect 14140 16258 14196 16268
rect 13804 16212 13860 16222
rect 13804 16118 13860 16156
rect 14364 16098 14420 16110
rect 14364 16046 14366 16098
rect 14418 16046 14420 16098
rect 13804 15876 13860 15886
rect 13468 15874 13860 15876
rect 13468 15822 13806 15874
rect 13858 15822 13860 15874
rect 13468 15820 13860 15822
rect 13804 15810 13860 15820
rect 13132 15204 13188 15214
rect 13132 15110 13188 15148
rect 14364 15204 14420 16046
rect 15036 15428 15092 16940
rect 16604 16098 16660 18396
rect 16940 18338 16996 19740
rect 16940 18286 16942 18338
rect 16994 18286 16996 18338
rect 16940 18274 16996 18286
rect 17052 18340 17108 20524
rect 18060 20018 18116 22428
rect 18060 19966 18062 20018
rect 18114 19966 18116 20018
rect 18060 19954 18116 19966
rect 18508 20018 18564 23548
rect 18732 22484 18788 22494
rect 18956 22484 19012 23662
rect 20188 23716 20244 23726
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20188 23268 20244 23660
rect 20188 23266 20692 23268
rect 20188 23214 20190 23266
rect 20242 23214 20692 23266
rect 20188 23212 20692 23214
rect 20188 23202 20244 23212
rect 18732 22482 19012 22484
rect 18732 22430 18734 22482
rect 18786 22430 19012 22482
rect 18732 22428 19012 22430
rect 19180 23154 19236 23166
rect 19180 23102 19182 23154
rect 19234 23102 19236 23154
rect 18732 22418 18788 22428
rect 18732 20690 18788 20702
rect 18732 20638 18734 20690
rect 18786 20638 18788 20690
rect 18732 20244 18788 20638
rect 18732 20178 18788 20188
rect 18508 19966 18510 20018
rect 18562 19966 18564 20018
rect 18508 19954 18564 19966
rect 18284 19908 18340 19918
rect 18284 19814 18340 19852
rect 17724 19794 17780 19806
rect 17724 19742 17726 19794
rect 17778 19742 17780 19794
rect 17052 18274 17108 18284
rect 17276 18340 17332 18350
rect 17276 17778 17332 18284
rect 17724 18228 17780 19742
rect 17836 19796 17892 19806
rect 17836 19702 17892 19740
rect 19180 19124 19236 23102
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20636 21812 20692 23212
rect 20860 22482 20916 25452
rect 20972 23716 21028 26910
rect 22316 26402 22372 27916
rect 22540 27906 22596 27916
rect 25004 27860 25060 27870
rect 25004 27766 25060 27804
rect 25564 27186 25620 28364
rect 25676 28084 25732 28590
rect 26124 28642 26180 28654
rect 26124 28590 26126 28642
rect 26178 28590 26180 28642
rect 25788 28420 25844 28430
rect 25788 28326 25844 28364
rect 25676 28028 25844 28084
rect 25676 27860 25732 27870
rect 25676 27766 25732 27804
rect 25564 27134 25566 27186
rect 25618 27134 25620 27186
rect 25564 27122 25620 27134
rect 24892 27074 24948 27086
rect 24892 27022 24894 27074
rect 24946 27022 24948 27074
rect 23212 26852 23268 26862
rect 22316 26350 22318 26402
rect 22370 26350 22372 26402
rect 22316 26338 22372 26350
rect 22988 26850 23268 26852
rect 22988 26798 23214 26850
rect 23266 26798 23268 26850
rect 22988 26796 23268 26798
rect 21644 26290 21700 26302
rect 21644 26238 21646 26290
rect 21698 26238 21700 26290
rect 21644 25508 21700 26238
rect 22988 25618 23044 26796
rect 23212 26786 23268 26796
rect 22988 25566 22990 25618
rect 23042 25566 23044 25618
rect 22988 25554 23044 25566
rect 23996 26516 24052 26526
rect 21644 25442 21700 25452
rect 22316 25508 22372 25518
rect 22316 25414 22372 25452
rect 23996 25508 24052 26460
rect 24892 26516 24948 27022
rect 24892 26384 24948 26460
rect 25564 26516 25620 26526
rect 24444 26180 24500 26190
rect 24444 26086 24500 26124
rect 25116 25620 25172 25630
rect 25116 25526 25172 25564
rect 25564 25618 25620 26460
rect 25564 25566 25566 25618
rect 25618 25566 25620 25618
rect 25564 25554 25620 25566
rect 25788 25620 25844 28028
rect 26124 26180 26180 28590
rect 26236 27972 26292 30718
rect 26572 30772 26628 30782
rect 26908 30772 26964 31838
rect 27020 30994 27076 32396
rect 27020 30942 27022 30994
rect 27074 30942 27076 30994
rect 27020 30930 27076 30942
rect 27356 31554 27412 31566
rect 27356 31502 27358 31554
rect 27410 31502 27412 31554
rect 26572 30770 26964 30772
rect 26572 30718 26574 30770
rect 26626 30718 26964 30770
rect 26572 30716 26964 30718
rect 26572 30706 26628 30716
rect 27244 29988 27300 29998
rect 27244 29538 27300 29932
rect 27244 29486 27246 29538
rect 27298 29486 27300 29538
rect 27244 29474 27300 29486
rect 26572 29428 26628 29438
rect 26572 29334 26628 29372
rect 27356 29428 27412 31502
rect 29708 30996 29764 32732
rect 32620 31948 32676 33406
rect 32508 31892 32676 31948
rect 32732 32676 32788 32686
rect 31948 31778 32004 31790
rect 31948 31726 31950 31778
rect 32002 31726 32004 31778
rect 31948 31556 32004 31726
rect 29708 30902 29764 30940
rect 29932 30996 29988 31006
rect 28140 29988 28196 29998
rect 28140 29894 28196 29932
rect 27356 29362 27412 29372
rect 28140 29428 28196 29438
rect 26348 28642 26404 28654
rect 26348 28590 26350 28642
rect 26402 28590 26404 28642
rect 26348 28084 26404 28590
rect 26348 28018 26404 28028
rect 27692 28084 27748 28094
rect 26236 27906 26292 27916
rect 26124 26114 26180 26124
rect 26348 27860 26404 27870
rect 25788 25554 25844 25564
rect 21756 24612 21812 24622
rect 21756 24518 21812 24556
rect 22204 24610 22260 24622
rect 22204 24558 22206 24610
rect 22258 24558 22260 24610
rect 20972 23650 21028 23660
rect 22204 23716 22260 24558
rect 23996 23938 24052 25452
rect 25676 24834 25732 24846
rect 25676 24782 25678 24834
rect 25730 24782 25732 24834
rect 24668 24052 24724 24062
rect 24668 23958 24724 23996
rect 25676 24052 25732 24782
rect 25676 23986 25732 23996
rect 23996 23886 23998 23938
rect 24050 23886 24052 23938
rect 23996 23874 24052 23886
rect 22204 23650 22260 23660
rect 26348 23378 26404 27804
rect 27692 27186 27748 28028
rect 27692 27134 27694 27186
rect 27746 27134 27748 27186
rect 27692 27122 27748 27134
rect 28140 26962 28196 29372
rect 29932 29426 29988 30940
rect 31948 30996 32004 31500
rect 32508 31556 32564 31892
rect 32620 31780 32676 31790
rect 32732 31780 32788 32620
rect 33628 32676 33684 32686
rect 33628 32582 33684 32620
rect 35868 32562 35924 34974
rect 36540 34690 36596 34702
rect 36540 34638 36542 34690
rect 36594 34638 36596 34690
rect 36540 34244 36596 34638
rect 36540 34178 36596 34188
rect 37436 34244 37492 34254
rect 37436 34150 37492 34188
rect 36428 34020 36484 34030
rect 36316 33346 36372 33358
rect 36316 33294 36318 33346
rect 36370 33294 36372 33346
rect 36316 33124 36372 33294
rect 36316 33058 36372 33068
rect 35868 32510 35870 32562
rect 35922 32510 35924 32562
rect 35868 32498 35924 32510
rect 36428 32562 36484 33964
rect 36540 33348 36596 33358
rect 36540 32674 36596 33292
rect 37660 33348 37716 37214
rect 37884 37266 37940 37884
rect 38332 37492 38388 37502
rect 38332 37398 38388 37436
rect 40684 37490 40740 37996
rect 41020 37986 41076 37996
rect 40684 37438 40686 37490
rect 40738 37438 40740 37490
rect 40684 37426 40740 37438
rect 41468 37490 41524 37996
rect 41468 37438 41470 37490
rect 41522 37438 41524 37490
rect 41468 37426 41524 37438
rect 37884 37214 37886 37266
rect 37938 37214 37940 37266
rect 37884 37202 37940 37214
rect 42364 37156 42420 37166
rect 42028 37154 42420 37156
rect 42028 37102 42366 37154
rect 42418 37102 42420 37154
rect 42028 37100 42420 37102
rect 39452 36482 39508 36494
rect 39452 36430 39454 36482
rect 39506 36430 39508 36482
rect 39452 35252 39508 36430
rect 40796 36484 40852 36494
rect 40124 36372 40180 36382
rect 40124 36370 40404 36372
rect 40124 36318 40126 36370
rect 40178 36318 40404 36370
rect 40124 36316 40404 36318
rect 40124 36306 40180 36316
rect 40348 35922 40404 36316
rect 40348 35870 40350 35922
rect 40402 35870 40404 35922
rect 40348 35858 40404 35870
rect 37996 34914 38052 34926
rect 37996 34862 37998 34914
rect 38050 34862 38052 34914
rect 37996 34132 38052 34862
rect 38668 34804 38724 34814
rect 38668 34802 38948 34804
rect 38668 34750 38670 34802
rect 38722 34750 38948 34802
rect 38668 34748 38948 34750
rect 38668 34738 38724 34748
rect 38892 34354 38948 34748
rect 38892 34302 38894 34354
rect 38946 34302 38948 34354
rect 38892 34290 38948 34302
rect 39452 34354 39508 35196
rect 39452 34302 39454 34354
rect 39506 34302 39508 34354
rect 38220 34132 38276 34142
rect 37996 34076 38220 34132
rect 38220 34038 38276 34076
rect 39452 34132 39508 34302
rect 39452 34066 39508 34076
rect 40572 35252 40628 35262
rect 37660 33282 37716 33292
rect 40572 33684 40628 35196
rect 40796 35026 40852 36428
rect 42028 36036 42084 37100
rect 42364 37090 42420 37100
rect 42812 37154 42868 38668
rect 42924 37492 42980 38782
rect 42924 37426 42980 37436
rect 43036 38834 43204 38836
rect 43036 38782 43150 38834
rect 43202 38782 43204 38834
rect 43036 38780 43204 38782
rect 42812 37102 42814 37154
rect 42866 37102 42868 37154
rect 42812 37090 42868 37102
rect 42252 36594 42308 36606
rect 42252 36542 42254 36594
rect 42306 36542 42308 36594
rect 42252 36484 42308 36542
rect 42924 36484 42980 36494
rect 42252 36482 42980 36484
rect 42252 36430 42926 36482
rect 42978 36430 42980 36482
rect 42252 36428 42980 36430
rect 42924 36418 42980 36428
rect 43036 36258 43092 38780
rect 43148 38770 43204 38780
rect 43484 38836 43540 38846
rect 43484 38742 43540 38780
rect 43932 38834 43988 38846
rect 43932 38782 43934 38834
rect 43986 38782 43988 38834
rect 43932 38162 43988 38782
rect 44156 38834 44212 39676
rect 44156 38782 44158 38834
rect 44210 38782 44212 38834
rect 44156 38770 44212 38782
rect 44604 38834 44660 40236
rect 45612 40290 45892 40292
rect 45612 40238 45838 40290
rect 45890 40238 45892 40290
rect 45612 40236 45892 40238
rect 45612 39506 45668 40236
rect 45836 40226 45892 40236
rect 46620 39732 46676 40350
rect 46620 39666 46676 39676
rect 45612 39454 45614 39506
rect 45666 39454 45668 39506
rect 45612 39442 45668 39454
rect 46844 39620 46900 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 49532 40402 49588 40414
rect 49532 40350 49534 40402
rect 49586 40350 49588 40402
rect 47628 39732 47684 39742
rect 47628 39638 47684 39676
rect 44604 38782 44606 38834
rect 44658 38782 44660 38834
rect 44604 38770 44660 38782
rect 46844 39394 46900 39564
rect 46844 39342 46846 39394
rect 46898 39342 46900 39394
rect 44380 38724 44436 38734
rect 44380 38630 44436 38668
rect 43932 38110 43934 38162
rect 43986 38110 43988 38162
rect 43932 38098 43988 38110
rect 44604 37828 44660 37838
rect 44604 37826 44996 37828
rect 44604 37774 44606 37826
rect 44658 37774 44996 37826
rect 44604 37772 44996 37774
rect 44604 37762 44660 37772
rect 44940 37378 44996 37772
rect 44940 37326 44942 37378
rect 44994 37326 44996 37378
rect 44940 37314 44996 37326
rect 45612 37268 45668 37278
rect 45500 37266 45668 37268
rect 45500 37214 45614 37266
rect 45666 37214 45668 37266
rect 45500 37212 45668 37214
rect 43484 36596 43540 36606
rect 43148 36484 43204 36494
rect 43148 36390 43204 36428
rect 43372 36482 43428 36494
rect 43372 36430 43374 36482
rect 43426 36430 43428 36482
rect 43036 36206 43038 36258
rect 43090 36206 43092 36258
rect 43036 36194 43092 36206
rect 41468 35980 42084 36036
rect 41468 35922 41524 35980
rect 41468 35870 41470 35922
rect 41522 35870 41524 35922
rect 41468 35252 41524 35870
rect 41468 35186 41524 35196
rect 41804 35364 41860 35374
rect 40796 34974 40798 35026
rect 40850 34974 40852 35026
rect 40796 34962 40852 34974
rect 41804 35026 41860 35308
rect 41804 34974 41806 35026
rect 41858 34974 41860 35026
rect 41804 34962 41860 34974
rect 41356 34690 41412 34702
rect 41356 34638 41358 34690
rect 41410 34638 41412 34690
rect 40796 34244 40852 34254
rect 40796 34242 41300 34244
rect 40796 34190 40798 34242
rect 40850 34190 41300 34242
rect 40796 34188 41300 34190
rect 40796 34178 40852 34188
rect 40572 33346 40628 33628
rect 41244 33458 41300 34188
rect 41244 33406 41246 33458
rect 41298 33406 41300 33458
rect 41244 33394 41300 33406
rect 41356 34132 41412 34638
rect 40572 33294 40574 33346
rect 40626 33294 40628 33346
rect 40572 33282 40628 33294
rect 36764 33124 36820 33134
rect 36764 33030 36820 33068
rect 37660 33124 37716 33134
rect 36540 32622 36542 32674
rect 36594 32622 36596 32674
rect 36540 32610 36596 32622
rect 36428 32510 36430 32562
rect 36482 32510 36484 32562
rect 36428 32498 36484 32510
rect 34748 32340 34804 32350
rect 34748 31890 34804 32284
rect 35980 32340 36036 32350
rect 35980 32246 36036 32284
rect 36204 32338 36260 32350
rect 36204 32286 36206 32338
rect 36258 32286 36260 32338
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 36204 31948 36260 32286
rect 36204 31892 36596 31948
rect 34748 31838 34750 31890
rect 34802 31838 34804 31890
rect 34748 31826 34804 31838
rect 32620 31778 32788 31780
rect 32620 31726 32622 31778
rect 32674 31726 32788 31778
rect 32620 31724 32788 31726
rect 32620 31714 32676 31724
rect 32508 31490 32564 31500
rect 33740 31556 33796 31566
rect 33740 30996 33796 31500
rect 35196 31556 35252 31566
rect 35196 31462 35252 31500
rect 31948 30930 32004 30940
rect 33292 30994 33796 30996
rect 33292 30942 33742 30994
rect 33794 30942 33796 30994
rect 33292 30940 33796 30942
rect 30380 30884 30436 30894
rect 30044 30882 30436 30884
rect 30044 30830 30382 30882
rect 30434 30830 30436 30882
rect 30044 30828 30436 30830
rect 30044 30098 30100 30828
rect 30380 30818 30436 30828
rect 32508 30882 32564 30894
rect 32508 30830 32510 30882
rect 32562 30830 32564 30882
rect 32284 30324 32340 30334
rect 32284 30230 32340 30268
rect 30044 30046 30046 30098
rect 30098 30046 30100 30098
rect 30044 30034 30100 30046
rect 29932 29374 29934 29426
rect 29986 29374 29988 29426
rect 29932 29362 29988 29374
rect 30492 29986 30548 29998
rect 31724 29988 31780 29998
rect 30492 29934 30494 29986
rect 30546 29934 30548 29986
rect 29372 29314 29428 29326
rect 29372 29262 29374 29314
rect 29426 29262 29428 29314
rect 28252 28644 28308 28654
rect 28252 28550 28308 28588
rect 28812 28420 28868 28430
rect 28812 28418 29316 28420
rect 28812 28366 28814 28418
rect 28866 28366 29316 28418
rect 28812 28364 29316 28366
rect 28812 28354 28868 28364
rect 28140 26910 28142 26962
rect 28194 26910 28196 26962
rect 28140 26516 28196 26910
rect 28028 26460 28140 26516
rect 27468 24722 27524 24734
rect 27468 24670 27470 24722
rect 27522 24670 27524 24722
rect 26796 24052 26852 24062
rect 26796 23958 26852 23996
rect 26348 23326 26350 23378
rect 26402 23326 26404 23378
rect 20860 22430 20862 22482
rect 20914 22430 20916 22482
rect 20860 22418 20916 22430
rect 23436 23268 23492 23278
rect 21644 22370 21700 22382
rect 21644 22318 21646 22370
rect 21698 22318 21700 22370
rect 20860 21812 20916 21822
rect 21308 21812 21364 21822
rect 21644 21812 21700 22318
rect 22428 22258 22484 22270
rect 22428 22206 22430 22258
rect 22482 22206 22484 22258
rect 20636 21810 21700 21812
rect 20636 21758 20862 21810
rect 20914 21758 21310 21810
rect 21362 21758 21700 21810
rect 20636 21756 21700 21758
rect 22316 21812 22372 21822
rect 22428 21812 22484 22206
rect 22316 21810 22484 21812
rect 22316 21758 22318 21810
rect 22370 21758 22484 21810
rect 22316 21756 22484 21758
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19516 20244 19572 20254
rect 19516 20150 19572 20188
rect 20636 20242 20692 21756
rect 20860 21746 20916 21756
rect 21308 21746 21364 21756
rect 22316 21746 22372 21756
rect 23212 21700 23268 21710
rect 20860 20916 20916 20926
rect 20860 20822 20916 20860
rect 23212 20914 23268 21644
rect 23212 20862 23214 20914
rect 23266 20862 23268 20914
rect 23212 20850 23268 20862
rect 22540 20802 22596 20814
rect 22540 20750 22542 20802
rect 22594 20750 22596 20802
rect 20636 20190 20638 20242
rect 20690 20190 20692 20242
rect 20636 20178 20692 20190
rect 21868 20578 21924 20590
rect 21868 20526 21870 20578
rect 21922 20526 21924 20578
rect 21868 20132 21924 20526
rect 21980 20132 22036 20142
rect 21868 20130 22036 20132
rect 21868 20078 21982 20130
rect 22034 20078 22036 20130
rect 21868 20076 22036 20078
rect 21980 20066 22036 20076
rect 21196 20018 21252 20030
rect 21196 19966 21198 20018
rect 21250 19966 21252 20018
rect 19180 19058 19236 19068
rect 19516 19124 19572 19134
rect 19404 18564 19460 18574
rect 17948 18452 18004 18462
rect 17948 18358 18004 18396
rect 18620 18340 18676 18350
rect 18620 18338 18900 18340
rect 18620 18286 18622 18338
rect 18674 18286 18900 18338
rect 18620 18284 18900 18286
rect 18620 18274 18676 18284
rect 17724 18162 17780 18172
rect 17276 17726 17278 17778
rect 17330 17726 17332 17778
rect 17276 17714 17332 17726
rect 18844 17554 18900 18284
rect 18844 17502 18846 17554
rect 18898 17502 18900 17554
rect 18844 17490 18900 17502
rect 17724 16996 17780 17006
rect 17276 16994 17780 16996
rect 17276 16942 17726 16994
rect 17778 16942 17780 16994
rect 17276 16940 17780 16942
rect 17276 16210 17332 16940
rect 17724 16930 17780 16940
rect 17276 16158 17278 16210
rect 17330 16158 17332 16210
rect 17276 16146 17332 16158
rect 19292 16884 19348 16894
rect 19292 16212 19348 16828
rect 19404 16882 19460 18508
rect 19404 16830 19406 16882
rect 19458 16830 19460 16882
rect 19404 16818 19460 16830
rect 19516 17892 19572 19068
rect 20076 19124 20132 19134
rect 20076 19030 20132 19068
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 21196 18564 21252 19966
rect 22540 19908 22596 20750
rect 21532 19348 21588 19358
rect 21532 19254 21588 19292
rect 21196 18498 21252 18508
rect 22540 18564 22596 19852
rect 22988 19348 23044 19358
rect 23436 19348 23492 23212
rect 26348 23268 26404 23326
rect 26348 23202 26404 23212
rect 26684 23716 26740 23726
rect 24556 22484 24612 22494
rect 24108 22482 24612 22484
rect 24108 22430 24558 22482
rect 24610 22430 24612 22482
rect 24108 22428 24612 22430
rect 23996 21812 24052 21822
rect 22988 19346 23492 19348
rect 22988 19294 22990 19346
rect 23042 19294 23492 19346
rect 22988 19292 23492 19294
rect 22988 19124 23044 19292
rect 23436 19236 23492 19292
rect 23660 21810 24052 21812
rect 23660 21758 23998 21810
rect 24050 21758 24052 21810
rect 23660 21756 24052 21758
rect 23548 19236 23604 19246
rect 23436 19234 23604 19236
rect 23436 19182 23550 19234
rect 23602 19182 23604 19234
rect 23436 19180 23604 19182
rect 23548 19170 23604 19180
rect 22988 19058 23044 19068
rect 23660 19012 23716 21756
rect 23996 21746 24052 21756
rect 24108 21586 24164 22428
rect 24556 22418 24612 22428
rect 26684 22482 26740 23660
rect 27356 23716 27412 23726
rect 27356 23622 27412 23660
rect 26908 23156 26964 23166
rect 26684 22430 26686 22482
rect 26738 22430 26740 22482
rect 26684 22418 26740 22430
rect 26796 23100 26908 23156
rect 26012 22372 26068 22382
rect 25676 21700 25732 21710
rect 25676 21606 25732 21644
rect 24108 21534 24110 21586
rect 24162 21534 24164 21586
rect 24108 21522 24164 21534
rect 23996 21362 24052 21374
rect 23996 21310 23998 21362
rect 24050 21310 24052 21362
rect 23996 19908 24052 21310
rect 24332 21362 24388 21374
rect 24332 21310 24334 21362
rect 24386 21310 24388 21362
rect 24332 20916 24388 21310
rect 24332 20850 24388 20860
rect 24556 21362 24612 21374
rect 24556 21310 24558 21362
rect 24610 21310 24612 21362
rect 24556 20916 24612 21310
rect 24556 20850 24612 20860
rect 25340 20916 25396 20926
rect 25340 20822 25396 20860
rect 26012 20802 26068 22316
rect 26012 20750 26014 20802
rect 26066 20750 26068 20802
rect 26012 20738 26068 20750
rect 26684 20690 26740 20702
rect 26684 20638 26686 20690
rect 26738 20638 26740 20690
rect 26684 20244 26740 20638
rect 26684 20178 26740 20188
rect 24108 19908 24164 19918
rect 23996 19906 24164 19908
rect 23996 19854 24110 19906
rect 24162 19854 24164 19906
rect 23996 19852 24164 19854
rect 24108 19842 24164 19852
rect 24556 19908 24612 19918
rect 24556 19814 24612 19852
rect 25452 19908 25508 19918
rect 25564 19908 25620 19918
rect 25508 19906 25620 19908
rect 25508 19854 25566 19906
rect 25618 19854 25620 19906
rect 25508 19852 25620 19854
rect 23548 18956 23716 19012
rect 25452 19124 25508 19852
rect 25564 19842 25620 19852
rect 25564 19124 25620 19134
rect 25452 19122 25620 19124
rect 25452 19070 25566 19122
rect 25618 19070 25620 19122
rect 25452 19068 25620 19070
rect 22540 18498 22596 18508
rect 22764 18564 22820 18574
rect 19404 16212 19460 16222
rect 19292 16210 19460 16212
rect 19292 16158 19406 16210
rect 19458 16158 19460 16210
rect 19292 16156 19460 16158
rect 19404 16146 19460 16156
rect 16604 16046 16606 16098
rect 16658 16046 16660 16098
rect 16604 16034 16660 16046
rect 15260 15428 15316 15438
rect 15036 15426 15316 15428
rect 15036 15374 15262 15426
rect 15314 15374 15316 15426
rect 15036 15372 15316 15374
rect 15260 15362 15316 15372
rect 14364 15138 14420 15148
rect 16044 15314 16100 15326
rect 16044 15262 16046 15314
rect 16098 15262 16100 15314
rect 16044 14308 16100 15262
rect 18844 15316 18900 15326
rect 18844 15222 18900 15260
rect 19516 15316 19572 17836
rect 19628 18452 19684 18462
rect 19628 16772 19684 18396
rect 21308 18452 21364 18462
rect 21308 18358 21364 18396
rect 21756 18450 21812 18462
rect 21756 18398 21758 18450
rect 21810 18398 21812 18450
rect 20748 18340 20804 18350
rect 20748 18246 20804 18284
rect 20188 17442 20244 17454
rect 20188 17390 20190 17442
rect 20242 17390 20244 17442
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20076 16996 20132 17006
rect 20188 16996 20244 17390
rect 20076 16994 20244 16996
rect 20076 16942 20078 16994
rect 20130 16942 20244 16994
rect 20076 16940 20244 16942
rect 20076 16930 20132 16940
rect 21756 16884 21812 18398
rect 21980 18340 22036 18350
rect 21980 18246 22036 18284
rect 21756 16818 21812 16828
rect 22204 18226 22260 18238
rect 22204 18174 22206 18226
rect 22258 18174 22260 18226
rect 19628 16716 19908 16772
rect 19852 16212 19908 16716
rect 22204 16770 22260 18174
rect 22428 18226 22484 18238
rect 22428 18174 22430 18226
rect 22482 18174 22484 18226
rect 22428 18004 22484 18174
rect 22540 18228 22596 18238
rect 22540 18134 22596 18172
rect 22428 17948 22708 18004
rect 22652 17778 22708 17948
rect 22652 17726 22654 17778
rect 22706 17726 22708 17778
rect 22652 17714 22708 17726
rect 22652 17108 22708 17118
rect 22764 17108 22820 18508
rect 22652 17106 22820 17108
rect 22652 17054 22654 17106
rect 22706 17054 22820 17106
rect 22652 17052 22820 17054
rect 23324 18228 23380 18238
rect 22652 17042 22708 17052
rect 23324 16882 23380 18172
rect 23324 16830 23326 16882
rect 23378 16830 23380 16882
rect 23324 16818 23380 16830
rect 22204 16718 22206 16770
rect 22258 16718 22260 16770
rect 22204 16706 22260 16718
rect 23548 16770 23604 18956
rect 23660 18564 23716 18574
rect 23660 18562 24836 18564
rect 23660 18510 23662 18562
rect 23714 18510 24836 18562
rect 23660 18508 24836 18510
rect 23660 18498 23716 18508
rect 24780 17778 24836 18508
rect 24780 17726 24782 17778
rect 24834 17726 24836 17778
rect 24780 17714 24836 17726
rect 25452 18452 25508 19068
rect 25564 19058 25620 19068
rect 25676 18452 25732 18462
rect 25452 18450 25732 18452
rect 25452 18398 25678 18450
rect 25730 18398 25732 18450
rect 25452 18396 25732 18398
rect 25452 17668 25508 18396
rect 25676 18386 25732 18396
rect 26460 18338 26516 18350
rect 26460 18286 26462 18338
rect 26514 18286 26516 18338
rect 25452 17666 25844 17668
rect 25452 17614 25454 17666
rect 25506 17614 25844 17666
rect 25452 17612 25844 17614
rect 25452 17602 25508 17612
rect 25788 17108 25844 17612
rect 26460 17554 26516 18286
rect 26460 17502 26462 17554
rect 26514 17502 26516 17554
rect 26460 17490 26516 17502
rect 25788 16976 25844 17052
rect 23548 16718 23550 16770
rect 23602 16718 23604 16770
rect 23548 16706 23604 16718
rect 23884 16658 23940 16670
rect 23884 16606 23886 16658
rect 23938 16606 23940 16658
rect 19852 16210 20244 16212
rect 19852 16158 19854 16210
rect 19906 16158 20244 16210
rect 19852 16156 20244 16158
rect 19852 16146 19908 16156
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 16604 15202 16660 15214
rect 16604 15150 16606 15202
rect 16658 15150 16660 15202
rect 19516 15184 19572 15260
rect 16604 14532 16660 15150
rect 20188 15092 20244 16156
rect 22540 15876 22596 15886
rect 19740 14644 19796 14654
rect 19516 14642 19796 14644
rect 19516 14590 19742 14642
rect 19794 14590 19796 14642
rect 19516 14588 19796 14590
rect 16828 14532 16884 14542
rect 16604 14530 16884 14532
rect 16604 14478 16830 14530
rect 16882 14478 16884 14530
rect 16604 14476 16884 14478
rect 16268 14308 16324 14318
rect 16044 14252 16268 14308
rect 16268 14214 16324 14252
rect 16828 14308 16884 14476
rect 17612 14420 17668 14430
rect 17612 14418 17892 14420
rect 17612 14366 17614 14418
rect 17666 14366 17892 14418
rect 17612 14364 17892 14366
rect 17612 14354 17668 14364
rect 16828 14242 16884 14252
rect 17276 14308 17332 14318
rect 12572 13682 12628 13692
rect 14028 13746 14084 13758
rect 14028 13694 14030 13746
rect 14082 13694 14084 13746
rect 11116 13634 11172 13646
rect 11116 13582 11118 13634
rect 11170 13582 11172 13634
rect 10668 12964 10724 12974
rect 11004 12964 11060 12974
rect 10668 12870 10724 12908
rect 10780 12962 11060 12964
rect 10780 12910 11006 12962
rect 11058 12910 11060 12962
rect 10780 12908 11060 12910
rect 10332 12290 10388 12796
rect 10332 12238 10334 12290
rect 10386 12238 10388 12290
rect 10332 12226 10388 12238
rect 9996 11564 10276 11620
rect 9996 11396 10052 11564
rect 9884 11394 10052 11396
rect 9884 11342 9998 11394
rect 10050 11342 10052 11394
rect 9884 11340 10052 11342
rect 9212 11172 9268 11182
rect 8988 11170 9268 11172
rect 8988 11118 9214 11170
rect 9266 11118 9268 11170
rect 8988 11116 9268 11118
rect 8596 9772 8708 9828
rect 8316 9716 8372 9726
rect 8316 9622 8372 9660
rect 8204 9214 8206 9266
rect 8258 9214 8260 9266
rect 8204 9202 8260 9214
rect 7644 9156 7700 9166
rect 7644 9062 7700 9100
rect 7196 8990 7198 9042
rect 7250 8990 7252 9042
rect 7196 8978 7252 8990
rect 7420 9044 7476 9054
rect 7420 8950 7476 8988
rect 7980 9044 8036 9054
rect 7980 8950 8036 8988
rect 8540 9044 8596 9772
rect 8652 9604 8708 9614
rect 8652 9154 8708 9548
rect 8652 9102 8654 9154
rect 8706 9102 8708 9154
rect 8652 9090 8708 9102
rect 8876 9156 8932 9166
rect 8540 8978 8596 8988
rect 8876 8428 8932 9100
rect 8988 8820 9044 8830
rect 8988 8726 9044 8764
rect 4956 8318 4958 8370
rect 5010 8318 5012 8370
rect 4956 8306 5012 8318
rect 6524 8372 6580 8382
rect 6524 8278 6580 8316
rect 8652 8372 8932 8428
rect 8652 8370 8708 8372
rect 8652 8318 8654 8370
rect 8706 8318 8708 8370
rect 8652 8306 8708 8318
rect 5740 8258 5796 8270
rect 5740 8206 5742 8258
rect 5794 8206 5796 8258
rect 3164 7534 3166 7586
rect 3218 7534 3220 7586
rect 3164 7522 3220 7534
rect 3948 7588 4004 7598
rect 3948 7494 4004 7532
rect 4844 7588 4900 7598
rect 2492 7420 2604 7476
rect 2604 7382 2660 7420
rect 2716 7474 2996 7476
rect 2716 7422 2830 7474
rect 2882 7422 2996 7474
rect 2716 7420 2996 7422
rect 3724 7476 3780 7486
rect 2268 6692 2324 6702
rect 2268 6598 2324 6636
rect 2716 6692 2772 7420
rect 2828 7410 2884 7420
rect 2716 6598 2772 6636
rect 3724 6580 3780 7420
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4172 6692 4228 6702
rect 4172 6598 4228 6636
rect 3724 6486 3780 6524
rect 2828 6466 2884 6478
rect 2828 6414 2830 6466
rect 2882 6414 2884 6466
rect 2828 6020 2884 6414
rect 2828 5954 2884 5964
rect 3948 6020 4004 6030
rect 3948 5926 4004 5964
rect 4732 5908 4788 5918
rect 4844 5908 4900 7532
rect 5740 7588 5796 8206
rect 9212 8036 9268 11116
rect 9772 10610 9828 10622
rect 9772 10558 9774 10610
rect 9826 10558 9828 10610
rect 9772 10500 9828 10558
rect 9772 10434 9828 10444
rect 9884 10164 9940 11340
rect 9996 11330 10052 11340
rect 10220 11396 10276 11406
rect 10220 11282 10276 11340
rect 10220 11230 10222 11282
rect 10274 11230 10276 11282
rect 10220 11218 10276 11230
rect 10668 11172 10724 11182
rect 10668 11078 10724 11116
rect 10780 10948 10836 12908
rect 11004 12898 11060 12908
rect 11004 12740 11060 12750
rect 11004 12646 11060 12684
rect 11004 12180 11060 12190
rect 11004 12086 11060 12124
rect 11116 11956 11172 13582
rect 12572 12964 12628 12974
rect 12572 12870 12628 12908
rect 12796 12962 12852 12974
rect 12796 12910 12798 12962
rect 12850 12910 12852 12962
rect 11340 12852 11396 12862
rect 11340 12758 11396 12796
rect 11900 12852 11956 12862
rect 11900 12758 11956 12796
rect 11676 12740 11732 12750
rect 11676 12290 11732 12684
rect 11676 12238 11678 12290
rect 11730 12238 11732 12290
rect 11676 12226 11732 12238
rect 11116 11890 11172 11900
rect 12124 11844 12180 11854
rect 11004 11172 11060 11182
rect 10108 10892 10948 10948
rect 10108 10834 10164 10892
rect 10108 10782 10110 10834
rect 10162 10782 10164 10834
rect 10108 10770 10164 10782
rect 10668 10722 10724 10734
rect 10668 10670 10670 10722
rect 10722 10670 10724 10722
rect 9884 9828 9940 10108
rect 9772 9826 9940 9828
rect 9772 9774 9886 9826
rect 9938 9774 9940 9826
rect 9772 9772 9940 9774
rect 8988 8034 9268 8036
rect 8988 7982 9214 8034
rect 9266 7982 9268 8034
rect 8988 7980 9268 7982
rect 5740 7522 5796 7532
rect 8540 7588 8596 7598
rect 8540 6690 8596 7532
rect 8988 7474 9044 7980
rect 9212 7970 9268 7980
rect 9324 9604 9380 9614
rect 9324 8260 9380 9548
rect 9772 9154 9828 9772
rect 9884 9762 9940 9772
rect 9996 10500 10052 10510
rect 9772 9102 9774 9154
rect 9826 9102 9828 9154
rect 9772 9090 9828 9102
rect 9996 9154 10052 10444
rect 10220 9604 10276 9614
rect 10220 9510 10276 9548
rect 9996 9102 9998 9154
rect 10050 9102 10052 9154
rect 9996 9090 10052 9102
rect 10108 9266 10164 9278
rect 10108 9214 10110 9266
rect 10162 9214 10164 9266
rect 10108 8372 10164 9214
rect 10556 9044 10612 9054
rect 10668 9044 10724 10670
rect 10892 9828 10948 10892
rect 11004 10612 11060 11116
rect 11900 11172 11956 11182
rect 11900 11078 11956 11116
rect 11004 10518 11060 10556
rect 12124 10722 12180 11788
rect 12796 11618 12852 12910
rect 13804 12964 13860 12974
rect 13356 12740 13412 12750
rect 13356 12180 13412 12684
rect 12796 11566 12798 11618
rect 12850 11566 12852 11618
rect 12796 11554 12852 11566
rect 13020 11844 13076 11854
rect 13020 11394 13076 11788
rect 13020 11342 13022 11394
rect 13074 11342 13076 11394
rect 13020 11330 13076 11342
rect 12236 11172 12292 11182
rect 12236 10834 12292 11116
rect 12460 11172 12516 11182
rect 12684 11172 12740 11182
rect 12460 11170 12628 11172
rect 12460 11118 12462 11170
rect 12514 11118 12628 11170
rect 12460 11116 12628 11118
rect 12460 11106 12516 11116
rect 12236 10782 12238 10834
rect 12290 10782 12292 10834
rect 12236 10770 12292 10782
rect 12124 10670 12126 10722
rect 12178 10670 12180 10722
rect 11228 10164 11284 10174
rect 11004 9828 11060 9838
rect 10892 9826 11172 9828
rect 10892 9774 11006 9826
rect 11058 9774 11172 9826
rect 10892 9772 11172 9774
rect 11004 9762 11060 9772
rect 10780 9714 10836 9726
rect 10780 9662 10782 9714
rect 10834 9662 10836 9714
rect 10780 9604 10836 9662
rect 10780 9268 10836 9548
rect 11004 9602 11060 9614
rect 11004 9550 11006 9602
rect 11058 9550 11060 9602
rect 10780 9212 10948 9268
rect 10556 9042 10724 9044
rect 10556 8990 10558 9042
rect 10610 8990 10724 9042
rect 10556 8988 10724 8990
rect 10556 8978 10612 8988
rect 10220 8820 10276 8830
rect 10220 8726 10276 8764
rect 10668 8428 10724 8988
rect 10892 8932 10948 9212
rect 11004 9156 11060 9550
rect 11004 9090 11060 9100
rect 11004 8932 11060 8942
rect 10892 8930 11060 8932
rect 10892 8878 11006 8930
rect 11058 8878 11060 8930
rect 10892 8876 11060 8878
rect 11004 8866 11060 8876
rect 11116 8428 11172 9772
rect 10668 8372 10836 8428
rect 10108 8306 10164 8316
rect 9660 8260 9716 8270
rect 9324 8258 9716 8260
rect 9324 8206 9662 8258
rect 9714 8206 9716 8258
rect 9324 8204 9716 8206
rect 9324 7700 9380 8204
rect 9660 8194 9716 8204
rect 10220 8258 10276 8270
rect 10220 8206 10222 8258
rect 10274 8206 10276 8258
rect 10108 8148 10164 8158
rect 10108 8054 10164 8092
rect 8988 7422 8990 7474
rect 9042 7422 9044 7474
rect 8988 7410 9044 7422
rect 9100 7644 9380 7700
rect 9884 8034 9940 8046
rect 9884 7982 9886 8034
rect 9938 7982 9940 8034
rect 8540 6638 8542 6690
rect 8594 6638 8596 6690
rect 8540 6626 8596 6638
rect 9100 6580 9156 7644
rect 9884 7364 9940 7982
rect 9212 7308 9940 7364
rect 9212 6802 9268 7308
rect 10220 7250 10276 8206
rect 10780 7364 10836 8372
rect 11004 8372 11172 8428
rect 11228 8428 11284 10108
rect 11340 9716 11396 9726
rect 11340 9622 11396 9660
rect 11900 9716 11956 9726
rect 11900 9622 11956 9660
rect 12124 8428 12180 10670
rect 12236 10386 12292 10398
rect 12236 10334 12238 10386
rect 12290 10334 12292 10386
rect 12236 9938 12292 10334
rect 12236 9886 12238 9938
rect 12290 9886 12292 9938
rect 12236 9874 12292 9886
rect 12572 9828 12628 11116
rect 12740 11116 12852 11172
rect 12684 11078 12740 11116
rect 12796 10834 12852 11116
rect 12796 10782 12798 10834
rect 12850 10782 12852 10834
rect 12796 10770 12852 10782
rect 12572 9734 12628 9772
rect 12796 9044 12852 9054
rect 12796 8950 12852 8988
rect 13356 9044 13412 12124
rect 13804 12180 13860 12908
rect 14028 12740 14084 13694
rect 14812 13634 14868 13646
rect 14812 13582 14814 13634
rect 14866 13582 14868 13634
rect 14812 12852 14868 13582
rect 16940 13634 16996 13646
rect 16940 13582 16942 13634
rect 16994 13582 16996 13634
rect 16940 13188 16996 13582
rect 16940 13122 16996 13132
rect 14812 12786 14868 12796
rect 15596 12852 15652 12862
rect 15596 12758 15652 12796
rect 16716 12740 16772 12750
rect 14028 12646 14084 12684
rect 16492 12738 16772 12740
rect 16492 12686 16718 12738
rect 16770 12686 16772 12738
rect 16492 12684 16772 12686
rect 13804 12066 13860 12124
rect 13804 12014 13806 12066
rect 13858 12014 13860 12066
rect 13804 12002 13860 12014
rect 14364 12290 14420 12302
rect 14364 12238 14366 12290
rect 14418 12238 14420 12290
rect 14252 11956 14308 11966
rect 14252 11862 14308 11900
rect 14028 11172 14084 11182
rect 14028 11078 14084 11116
rect 14364 11172 14420 12238
rect 14476 12180 14532 12190
rect 14476 12086 14532 12124
rect 15260 12178 15316 12190
rect 15260 12126 15262 12178
rect 15314 12126 15316 12178
rect 14364 11106 14420 11116
rect 15260 10500 15316 12126
rect 15596 12178 15652 12190
rect 15596 12126 15598 12178
rect 15650 12126 15652 12178
rect 15596 11844 15652 12126
rect 15596 11778 15652 11788
rect 16156 11508 16212 11518
rect 16156 11394 16212 11452
rect 16156 11342 16158 11394
rect 16210 11342 16212 11394
rect 16156 11330 16212 11342
rect 15260 10444 15652 10500
rect 15596 9828 15652 10444
rect 16492 9938 16548 12684
rect 16716 12674 16772 12684
rect 17276 12738 17332 14252
rect 17836 13970 17892 14364
rect 17836 13918 17838 13970
rect 17890 13918 17892 13970
rect 17836 13906 17892 13918
rect 19292 13188 19348 13198
rect 19292 13094 19348 13132
rect 19516 13186 19572 14588
rect 19740 14578 19796 14588
rect 20188 14642 20244 15036
rect 20188 14590 20190 14642
rect 20242 14590 20244 14642
rect 20188 14578 20244 14590
rect 20412 15316 20468 15326
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19516 13134 19518 13186
rect 19570 13134 19572 13186
rect 19516 13122 19572 13134
rect 19068 13076 19124 13086
rect 17276 12686 17278 12738
rect 17330 12686 17332 12738
rect 16828 11284 16884 11294
rect 17276 11284 17332 12686
rect 16828 11282 17332 11284
rect 16828 11230 16830 11282
rect 16882 11230 17332 11282
rect 16828 11228 17332 11230
rect 18620 13074 19124 13076
rect 18620 13022 19070 13074
rect 19122 13022 19124 13074
rect 18620 13020 19124 13022
rect 16492 9886 16494 9938
rect 16546 9886 16548 9938
rect 16492 9874 16548 9886
rect 16716 10722 16772 10734
rect 16716 10670 16718 10722
rect 16770 10670 16772 10722
rect 13468 9156 13524 9166
rect 13468 9062 13524 9100
rect 13356 8978 13412 8988
rect 15484 9044 15540 9054
rect 11228 8372 11396 8428
rect 11004 8258 11060 8372
rect 11004 8206 11006 8258
rect 11058 8206 11060 8258
rect 11004 8148 11060 8206
rect 11340 8258 11396 8372
rect 11900 8372 12180 8428
rect 11340 8206 11342 8258
rect 11394 8206 11396 8258
rect 11340 8194 11396 8206
rect 11564 8260 11620 8270
rect 11788 8260 11844 8270
rect 11900 8260 11956 8372
rect 11564 8258 11732 8260
rect 11564 8206 11566 8258
rect 11618 8206 11732 8258
rect 11564 8204 11732 8206
rect 11564 8194 11620 8204
rect 11004 8082 11060 8092
rect 10892 7476 10948 7486
rect 10892 7474 11396 7476
rect 10892 7422 10894 7474
rect 10946 7422 11396 7474
rect 10892 7420 11396 7422
rect 10892 7410 10948 7420
rect 10780 7270 10836 7308
rect 10220 7198 10222 7250
rect 10274 7198 10276 7250
rect 10220 7186 10276 7198
rect 9212 6750 9214 6802
rect 9266 6750 9268 6802
rect 9212 6738 9268 6750
rect 11340 6804 11396 7420
rect 11340 6672 11396 6748
rect 11452 7364 11508 7374
rect 9100 6514 9156 6524
rect 4732 5906 4900 5908
rect 4732 5854 4734 5906
rect 4786 5854 4900 5906
rect 4732 5852 4900 5854
rect 11452 5906 11508 7308
rect 11676 6132 11732 8204
rect 11788 8258 11956 8260
rect 11788 8206 11790 8258
rect 11842 8206 11956 8258
rect 11788 8204 11956 8206
rect 11788 8194 11844 8204
rect 11900 6914 11956 8204
rect 12012 8146 12068 8158
rect 12012 8094 12014 8146
rect 12066 8094 12068 8146
rect 12012 7364 12068 8094
rect 12124 8034 12180 8046
rect 12124 7982 12126 8034
rect 12178 7982 12180 8034
rect 12124 7588 12180 7982
rect 12124 7522 12180 7532
rect 14700 7588 14756 7598
rect 14700 7494 14756 7532
rect 15484 7474 15540 8988
rect 15596 8930 15652 9772
rect 15708 9826 15764 9838
rect 15708 9774 15710 9826
rect 15762 9774 15764 9826
rect 15708 9044 15764 9774
rect 15708 8978 15764 8988
rect 16044 9044 16100 9054
rect 15596 8878 15598 8930
rect 15650 8878 15652 8930
rect 15596 8866 15652 8878
rect 16044 8428 16100 8988
rect 15932 8372 16100 8428
rect 16604 8372 16660 8382
rect 16716 8372 16772 10670
rect 16828 9940 16884 11228
rect 16828 9044 16884 9884
rect 18620 9938 18676 13020
rect 19068 13010 19124 13020
rect 19964 13076 20020 13086
rect 19964 12982 20020 13020
rect 18620 9886 18622 9938
rect 18674 9886 18676 9938
rect 18620 9874 18676 9886
rect 18844 12850 18900 12862
rect 18844 12798 18846 12850
rect 18898 12798 18900 12850
rect 16828 8978 16884 8988
rect 18844 8428 18900 12798
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19964 12180 20020 12190
rect 19068 12178 20020 12180
rect 19068 12126 19966 12178
rect 20018 12126 20020 12178
rect 19068 12124 20020 12126
rect 19068 10612 19124 12124
rect 19964 12114 20020 12124
rect 20412 11508 20468 15260
rect 21532 15202 21588 15214
rect 21532 15150 21534 15202
rect 21586 15150 21588 15202
rect 21532 15148 21588 15150
rect 20636 15092 20692 15102
rect 20636 13746 20692 15036
rect 21420 15092 21588 15148
rect 21756 15092 21812 15102
rect 21420 15026 21476 15036
rect 21756 14530 21812 15036
rect 22540 14642 22596 15820
rect 23772 15876 23828 15886
rect 23772 15782 23828 15820
rect 23884 15148 23940 16606
rect 26236 15314 26292 15326
rect 26236 15262 26238 15314
rect 26290 15262 26292 15314
rect 23884 15092 24388 15148
rect 22540 14590 22542 14642
rect 22594 14590 22596 14642
rect 22540 14578 22596 14590
rect 21756 14478 21758 14530
rect 21810 14478 21812 14530
rect 20860 14308 20916 14318
rect 20860 14306 21364 14308
rect 20860 14254 20862 14306
rect 20914 14254 21364 14306
rect 20860 14252 21364 14254
rect 20860 14242 20916 14252
rect 21308 13858 21364 14252
rect 21756 13972 21812 14478
rect 21756 13906 21812 13916
rect 23884 13972 23940 13982
rect 23884 13878 23940 13916
rect 21308 13806 21310 13858
rect 21362 13806 21364 13858
rect 21308 13794 21364 13806
rect 20636 13694 20638 13746
rect 20690 13694 20692 13746
rect 20636 13682 20692 13694
rect 23436 13634 23492 13646
rect 23436 13582 23438 13634
rect 23490 13582 23492 13634
rect 23324 13076 23380 13086
rect 23324 12982 23380 13020
rect 23212 12964 23268 12974
rect 22988 12962 23268 12964
rect 22988 12910 23214 12962
rect 23266 12910 23268 12962
rect 22988 12908 23268 12910
rect 23436 12964 23492 13582
rect 23548 12964 23604 12974
rect 23436 12962 23604 12964
rect 23436 12910 23550 12962
rect 23602 12910 23604 12962
rect 23436 12908 23604 12910
rect 21644 12740 21700 12750
rect 20748 12738 21700 12740
rect 20748 12686 21646 12738
rect 21698 12686 21700 12738
rect 20748 12684 21700 12686
rect 20748 12290 20804 12684
rect 21644 12674 21700 12684
rect 20748 12238 20750 12290
rect 20802 12238 20804 12290
rect 20748 12226 20804 12238
rect 22876 12068 22932 12078
rect 22988 12068 23044 12908
rect 23212 12898 23268 12908
rect 23548 12898 23604 12908
rect 23884 12738 23940 12750
rect 23884 12686 23886 12738
rect 23938 12686 23940 12738
rect 23884 12404 23940 12686
rect 24332 12404 24388 15092
rect 24668 14644 24724 14654
rect 24668 14550 24724 14588
rect 25340 14530 25396 14542
rect 25340 14478 25342 14530
rect 25394 14478 25396 14530
rect 25340 13524 25396 14478
rect 26012 14418 26068 14430
rect 26012 14366 26014 14418
rect 26066 14366 26068 14418
rect 26012 13970 26068 14366
rect 26012 13918 26014 13970
rect 26066 13918 26068 13970
rect 26012 13906 26068 13918
rect 25564 13524 25620 13534
rect 25340 13468 25564 13524
rect 23548 12402 23940 12404
rect 23548 12350 23886 12402
rect 23938 12350 23940 12402
rect 23548 12348 23940 12350
rect 23436 12068 23492 12078
rect 22876 12066 23044 12068
rect 22876 12014 22878 12066
rect 22930 12014 23044 12066
rect 22876 12012 23044 12014
rect 23324 12066 23492 12068
rect 23324 12014 23438 12066
rect 23490 12014 23492 12066
rect 23324 12012 23492 12014
rect 22876 12002 22932 12012
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19068 10610 19236 10612
rect 19068 10558 19070 10610
rect 19122 10558 19236 10610
rect 19068 10556 19236 10558
rect 19068 10546 19124 10556
rect 19068 9940 19124 9950
rect 19068 9846 19124 9884
rect 19068 9268 19124 9278
rect 19068 9174 19124 9212
rect 15484 7422 15486 7474
rect 15538 7422 15540 7474
rect 15484 7410 15540 7422
rect 15820 8258 15876 8270
rect 15820 8206 15822 8258
rect 15874 8206 15876 8258
rect 12572 7364 12628 7374
rect 12012 7298 12068 7308
rect 12460 7362 12628 7364
rect 12460 7310 12574 7362
rect 12626 7310 12628 7362
rect 12460 7308 12628 7310
rect 11900 6862 11902 6914
rect 11954 6862 11956 6914
rect 11900 6850 11956 6862
rect 12236 6804 12292 6814
rect 12236 6710 12292 6748
rect 11900 6692 11956 6702
rect 11788 6132 11844 6142
rect 11676 6130 11844 6132
rect 11676 6078 11790 6130
rect 11842 6078 11844 6130
rect 11676 6076 11844 6078
rect 11788 6066 11844 6076
rect 11900 6018 11956 6636
rect 12460 6690 12516 7308
rect 12572 7298 12628 7308
rect 12460 6638 12462 6690
rect 12514 6638 12516 6690
rect 11900 5966 11902 6018
rect 11954 5966 11956 6018
rect 11900 5954 11956 5966
rect 12124 6020 12180 6030
rect 12460 6020 12516 6638
rect 15820 6692 15876 8206
rect 15932 7698 15988 8372
rect 16604 8370 16772 8372
rect 16604 8318 16606 8370
rect 16658 8318 16772 8370
rect 16604 8316 16772 8318
rect 18732 8372 18900 8428
rect 18732 8370 18788 8372
rect 18732 8318 18734 8370
rect 18786 8318 18788 8370
rect 16604 8306 16660 8316
rect 18732 8306 18788 8318
rect 15932 7646 15934 7698
rect 15986 7646 15988 7698
rect 15932 7634 15988 7646
rect 19180 8034 19236 10556
rect 19740 10498 19796 10510
rect 19740 10446 19742 10498
rect 19794 10446 19796 10498
rect 19740 10276 19796 10446
rect 19740 10210 19796 10220
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20412 9268 20468 11452
rect 21980 11394 22036 11406
rect 21980 11342 21982 11394
rect 22034 11342 22036 11394
rect 21980 10612 22036 11342
rect 22316 11284 22372 11294
rect 22316 11282 22484 11284
rect 22316 11230 22318 11282
rect 22370 11230 22484 11282
rect 22316 11228 22484 11230
rect 22316 11218 22372 11228
rect 21868 10500 21924 10510
rect 21980 10500 22036 10556
rect 21868 10498 22036 10500
rect 21868 10446 21870 10498
rect 21922 10446 22036 10498
rect 21868 10444 22036 10446
rect 21868 10434 21924 10444
rect 20412 9042 20468 9212
rect 20412 8990 20414 9042
rect 20466 8990 20468 9042
rect 20412 8978 20468 8990
rect 21868 10276 21924 10286
rect 21756 8484 21812 8494
rect 21868 8484 21924 10220
rect 21980 9938 22036 10444
rect 22204 11170 22260 11182
rect 22204 11118 22206 11170
rect 22258 11118 22260 11170
rect 22204 10052 22260 11118
rect 22428 10610 22484 11228
rect 22876 10724 22932 10734
rect 22876 10722 23156 10724
rect 22876 10670 22878 10722
rect 22930 10670 23156 10722
rect 22876 10668 23156 10670
rect 22876 10658 22932 10668
rect 22428 10558 22430 10610
rect 22482 10558 22484 10610
rect 22204 9996 22372 10052
rect 21980 9886 21982 9938
rect 22034 9886 22036 9938
rect 21980 9874 22036 9886
rect 22204 9828 22260 9838
rect 22204 9734 22260 9772
rect 21756 8482 21924 8484
rect 21756 8430 21758 8482
rect 21810 8430 21924 8482
rect 21756 8428 21924 8430
rect 22092 8484 22148 8522
rect 21756 8418 21812 8428
rect 22092 8418 22148 8428
rect 20860 8260 20916 8270
rect 20860 8166 20916 8204
rect 21868 8260 21924 8270
rect 21868 8166 21924 8204
rect 22316 8258 22372 9996
rect 22428 9828 22484 10558
rect 22652 10612 22708 10622
rect 22652 10518 22708 10556
rect 22988 10500 23044 10510
rect 22988 10406 23044 10444
rect 22428 9762 22484 9772
rect 22540 9604 22596 9614
rect 22540 9602 22932 9604
rect 22540 9550 22542 9602
rect 22594 9550 22932 9602
rect 22540 9548 22932 9550
rect 22540 9538 22596 9548
rect 22876 8484 22932 9548
rect 22876 8418 22932 8428
rect 22316 8206 22318 8258
rect 22370 8206 22372 8258
rect 22316 8194 22372 8206
rect 19180 7982 19182 8034
rect 19234 7982 19236 8034
rect 15820 6626 15876 6636
rect 19180 7474 19236 7982
rect 19180 7422 19182 7474
rect 19234 7422 19236 7474
rect 19180 6692 19236 7422
rect 12124 6018 12516 6020
rect 12124 5966 12126 6018
rect 12178 5966 12516 6018
rect 12124 5964 12516 5966
rect 12124 5954 12180 5964
rect 11452 5854 11454 5906
rect 11506 5854 11508 5906
rect 4732 5842 4788 5852
rect 11452 5842 11508 5854
rect 19180 5906 19236 6636
rect 19628 8036 19684 8046
rect 19628 6020 19684 7980
rect 20636 8034 20692 8046
rect 20636 7982 20638 8034
rect 20690 7982 20692 8034
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20636 7476 20692 7982
rect 20748 8036 20804 8046
rect 20748 7942 20804 7980
rect 22988 8034 23044 8046
rect 22988 7982 22990 8034
rect 23042 7982 23044 8034
rect 22764 7586 22820 7598
rect 22764 7534 22766 7586
rect 22818 7534 22820 7586
rect 20636 7410 20692 7420
rect 22092 7476 22148 7486
rect 19964 7364 20020 7374
rect 19964 7270 20020 7308
rect 22092 7362 22148 7420
rect 22092 7310 22094 7362
rect 22146 7310 22148 7362
rect 22092 7298 22148 7310
rect 22652 7364 22708 7374
rect 22652 7270 22708 7308
rect 22764 7252 22820 7534
rect 22988 7586 23044 7982
rect 22988 7534 22990 7586
rect 23042 7534 23044 7586
rect 22988 7522 23044 7534
rect 23100 8034 23156 10668
rect 23324 10500 23380 12012
rect 23436 12002 23492 12012
rect 23548 11394 23604 12348
rect 23884 12338 23940 12348
rect 23996 12348 24388 12404
rect 23996 12180 24052 12348
rect 24332 12290 24388 12348
rect 24332 12238 24334 12290
rect 24386 12238 24388 12290
rect 24332 12226 24388 12238
rect 23548 11342 23550 11394
rect 23602 11342 23604 11394
rect 23548 11330 23604 11342
rect 23660 12124 24052 12180
rect 24108 12180 24164 12190
rect 23660 11282 23716 12124
rect 24108 11396 24164 12124
rect 24220 11956 24276 11966
rect 24220 11954 24500 11956
rect 24220 11902 24222 11954
rect 24274 11902 24500 11954
rect 24220 11900 24500 11902
rect 24220 11890 24276 11900
rect 24220 11396 24276 11406
rect 24108 11394 24276 11396
rect 24108 11342 24222 11394
rect 24274 11342 24276 11394
rect 24108 11340 24276 11342
rect 24220 11330 24276 11340
rect 23660 11230 23662 11282
rect 23714 11230 23716 11282
rect 23660 11218 23716 11230
rect 23100 7982 23102 8034
rect 23154 7982 23156 8034
rect 23100 7476 23156 7982
rect 23100 7410 23156 7420
rect 23212 10498 23380 10500
rect 23212 10446 23326 10498
rect 23378 10446 23380 10498
rect 23212 10444 23380 10446
rect 23212 8930 23268 10444
rect 23324 10434 23380 10444
rect 23212 8878 23214 8930
rect 23266 8878 23268 8930
rect 22652 6804 22708 6814
rect 22764 6804 22820 7196
rect 22652 6802 22820 6804
rect 22652 6750 22654 6802
rect 22706 6750 22820 6802
rect 22652 6748 22820 6750
rect 22652 6738 22708 6748
rect 22092 6692 22148 6702
rect 22092 6466 22148 6636
rect 22092 6414 22094 6466
rect 22146 6414 22148 6466
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 22092 6132 22148 6414
rect 23212 6690 23268 8878
rect 24444 10050 24500 11900
rect 25004 11620 25060 11630
rect 25004 11526 25060 11564
rect 25452 11620 25508 11630
rect 24668 11394 24724 11406
rect 24668 11342 24670 11394
rect 24722 11342 24724 11394
rect 24668 10500 24724 11342
rect 24668 10434 24724 10444
rect 24444 9998 24446 10050
rect 24498 9998 24500 10050
rect 23996 8258 24052 8270
rect 23996 8206 23998 8258
rect 24050 8206 24052 8258
rect 23212 6638 23214 6690
rect 23266 6638 23268 6690
rect 22092 6066 22148 6076
rect 22428 6132 22484 6142
rect 22428 6038 22484 6076
rect 23212 6132 23268 6638
rect 23212 6066 23268 6076
rect 23660 7364 23716 7374
rect 23996 7364 24052 8206
rect 24444 8260 24500 9998
rect 24668 9828 24724 9838
rect 24668 9268 24724 9772
rect 24892 9828 24948 9838
rect 24892 9734 24948 9772
rect 24668 9202 24724 9212
rect 24780 9602 24836 9614
rect 24780 9550 24782 9602
rect 24834 9550 24836 9602
rect 24780 8370 24836 9550
rect 25452 8428 25508 11564
rect 25564 11394 25620 13468
rect 26236 13524 26292 15262
rect 26796 14980 26852 23100
rect 26908 23062 26964 23100
rect 27468 23044 27524 24670
rect 28028 24050 28084 26460
rect 28140 26450 28196 26460
rect 28588 26516 28644 26526
rect 28588 26290 28644 26460
rect 29260 26402 29316 28364
rect 29372 27860 29428 29262
rect 30268 28644 30324 28654
rect 30268 28550 30324 28588
rect 29372 27794 29428 27804
rect 30492 27970 30548 29934
rect 30716 29986 31780 29988
rect 30716 29934 31726 29986
rect 31778 29934 31780 29986
rect 30716 29932 31780 29934
rect 30716 29538 30772 29932
rect 31724 29922 31780 29932
rect 32508 29652 32564 30830
rect 32732 30324 32788 30334
rect 32732 30230 32788 30268
rect 33292 30324 33348 30940
rect 33740 30930 33796 30940
rect 34412 30884 34468 30894
rect 33292 30192 33348 30268
rect 34076 30882 34468 30884
rect 34076 30830 34414 30882
rect 34466 30830 34468 30882
rect 34076 30828 34468 30830
rect 34076 30098 34132 30828
rect 34412 30818 34468 30828
rect 36540 30882 36596 31892
rect 37548 31778 37604 31790
rect 37548 31726 37550 31778
rect 37602 31726 37604 31778
rect 36764 31554 36820 31566
rect 36764 31502 36766 31554
rect 36818 31502 36820 31554
rect 36764 31108 36820 31502
rect 36764 31042 36820 31052
rect 37100 30996 37156 31006
rect 37548 30996 37604 31726
rect 36540 30830 36542 30882
rect 36594 30830 36596 30882
rect 36540 30818 36596 30830
rect 36988 30994 37604 30996
rect 36988 30942 37102 30994
rect 37154 30942 37604 30994
rect 36988 30940 37604 30942
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34076 30046 34078 30098
rect 34130 30046 34132 30098
rect 34076 30034 34132 30046
rect 36988 30100 37044 30940
rect 37100 30930 37156 30940
rect 37660 30212 37716 33068
rect 37996 32674 38052 32686
rect 37996 32622 37998 32674
rect 38050 32622 38052 32674
rect 37996 31948 38052 32622
rect 37996 31892 38388 31948
rect 40460 31892 40516 31902
rect 38332 31890 38388 31892
rect 38332 31838 38334 31890
rect 38386 31838 38388 31890
rect 38332 31826 38388 31838
rect 40236 31890 40516 31892
rect 40236 31838 40462 31890
rect 40514 31838 40516 31890
rect 40236 31836 40516 31838
rect 37884 31108 37940 31118
rect 37884 31014 37940 31052
rect 40012 30884 40068 30894
rect 39452 30882 40068 30884
rect 39452 30830 40014 30882
rect 40066 30830 40068 30882
rect 39452 30828 40068 30830
rect 37660 30146 37716 30156
rect 38556 30212 38612 30222
rect 38556 30118 38612 30156
rect 30716 29486 30718 29538
rect 30770 29486 30772 29538
rect 30716 29474 30772 29486
rect 32060 29596 32564 29652
rect 32060 28532 32116 29596
rect 33740 29428 33796 29438
rect 33740 29334 33796 29372
rect 36988 29428 37044 30044
rect 36988 29334 37044 29372
rect 39452 29426 39508 30828
rect 40012 30818 40068 30828
rect 39452 29374 39454 29426
rect 39506 29374 39508 29426
rect 39452 29362 39508 29374
rect 39676 30324 39732 30334
rect 39676 29426 39732 30268
rect 40236 30324 40292 31836
rect 40460 31826 40516 31836
rect 40908 31556 40964 31566
rect 40796 31554 40964 31556
rect 40796 31502 40910 31554
rect 40962 31502 40964 31554
rect 40796 31500 40964 31502
rect 40460 30884 40516 30894
rect 40236 30258 40292 30268
rect 40348 30882 40516 30884
rect 40348 30830 40462 30882
rect 40514 30830 40516 30882
rect 40348 30828 40516 30830
rect 40348 30100 40404 30828
rect 40460 30818 40516 30828
rect 40348 30006 40404 30044
rect 40796 30100 40852 31500
rect 40908 31490 40964 31500
rect 39676 29374 39678 29426
rect 39730 29374 39732 29426
rect 39676 29362 39732 29374
rect 40796 29650 40852 30044
rect 40796 29598 40798 29650
rect 40850 29598 40852 29650
rect 40796 29428 40852 29598
rect 40796 29362 40852 29372
rect 32844 29316 32900 29326
rect 30492 27918 30494 27970
rect 30546 27918 30548 27970
rect 30492 26516 30548 27918
rect 31724 28476 32116 28532
rect 32172 29314 32900 29316
rect 32172 29262 32846 29314
rect 32898 29262 32900 29314
rect 32172 29260 32900 29262
rect 31500 27860 31556 27870
rect 31500 27766 31556 27804
rect 31724 27858 31780 28476
rect 31724 27806 31726 27858
rect 31778 27806 31780 27858
rect 31724 27794 31780 27806
rect 32060 28082 32116 28094
rect 32060 28030 32062 28082
rect 32114 28030 32116 28082
rect 30492 26450 30548 26460
rect 31388 27636 31444 27646
rect 29260 26350 29262 26402
rect 29314 26350 29316 26402
rect 29260 26338 29316 26350
rect 28588 26238 28590 26290
rect 28642 26238 28644 26290
rect 28588 26226 28644 26238
rect 31388 26178 31444 27580
rect 31948 27636 32004 27646
rect 31948 27542 32004 27580
rect 31836 26516 31892 26526
rect 31836 26422 31892 26460
rect 31388 26126 31390 26178
rect 31442 26126 31444 26178
rect 31388 26114 31444 26126
rect 32060 25732 32116 28030
rect 32172 27858 32228 29260
rect 32844 29250 32900 29260
rect 34412 29314 34468 29326
rect 34412 29262 34414 29314
rect 34466 29262 34468 29314
rect 32172 27806 32174 27858
rect 32226 27806 32228 27858
rect 32172 27794 32228 27806
rect 33404 28756 33460 28766
rect 32284 27186 32340 27198
rect 32284 27134 32286 27186
rect 32338 27134 32340 27186
rect 32284 26964 32340 27134
rect 32284 26898 32340 26908
rect 32396 26404 32452 26414
rect 31724 25676 32116 25732
rect 32172 26402 32452 26404
rect 32172 26350 32398 26402
rect 32450 26350 32452 26402
rect 32172 26348 32452 26350
rect 31388 25508 31444 25518
rect 31276 25452 31388 25508
rect 28252 25282 28308 25294
rect 28252 25230 28254 25282
rect 28306 25230 28308 25282
rect 28140 24836 28196 24846
rect 28252 24836 28308 25230
rect 28140 24834 28308 24836
rect 28140 24782 28142 24834
rect 28194 24782 28308 24834
rect 28140 24780 28308 24782
rect 28140 24770 28196 24780
rect 30268 24612 30324 24622
rect 30044 24610 30324 24612
rect 30044 24558 30270 24610
rect 30322 24558 30324 24610
rect 30044 24556 30324 24558
rect 30044 24162 30100 24556
rect 30268 24546 30324 24556
rect 30044 24110 30046 24162
rect 30098 24110 30100 24162
rect 30044 24098 30100 24110
rect 28028 23998 28030 24050
rect 28082 23998 28084 24050
rect 28028 23986 28084 23998
rect 29708 24052 29764 24062
rect 29708 23958 29764 23996
rect 29820 23938 29876 23950
rect 29820 23886 29822 23938
rect 29874 23886 29876 23938
rect 28476 23714 28532 23726
rect 28476 23662 28478 23714
rect 28530 23662 28532 23714
rect 27692 23044 27748 23054
rect 27468 22988 27692 23044
rect 27692 22372 27748 22988
rect 27692 21586 27748 22316
rect 28364 21700 28420 21710
rect 28476 21700 28532 23662
rect 29820 23268 29876 23886
rect 28812 23212 29876 23268
rect 30268 23938 30324 23950
rect 30268 23886 30270 23938
rect 30322 23886 30324 23938
rect 28812 22482 28868 23212
rect 28924 23044 28980 23054
rect 28924 22950 28980 22988
rect 30268 22708 30324 23886
rect 30380 23828 30436 23838
rect 30380 23734 30436 23772
rect 30268 22652 30548 22708
rect 28812 22430 28814 22482
rect 28866 22430 28868 22482
rect 28812 22418 28868 22430
rect 28364 21698 28532 21700
rect 28364 21646 28366 21698
rect 28418 21646 28532 21698
rect 28364 21644 28532 21646
rect 28364 21634 28420 21644
rect 27692 21534 27694 21586
rect 27746 21534 27748 21586
rect 27692 21522 27748 21534
rect 30492 21474 30548 22652
rect 31164 22372 31220 22382
rect 31276 22372 31332 25452
rect 31388 25376 31444 25452
rect 31164 22370 31332 22372
rect 31164 22318 31166 22370
rect 31218 22318 31332 22370
rect 31164 22316 31332 22318
rect 31388 23938 31444 23950
rect 31388 23886 31390 23938
rect 31442 23886 31444 23938
rect 31164 22306 31220 22316
rect 30492 21422 30494 21474
rect 30546 21422 30548 21474
rect 30492 21410 30548 21422
rect 28812 20914 28868 20926
rect 28812 20862 28814 20914
rect 28866 20862 28868 20914
rect 27468 20244 27524 20282
rect 27468 20178 27524 20188
rect 28812 20020 28868 20862
rect 31164 20916 31220 20926
rect 29708 20802 29764 20814
rect 29708 20750 29710 20802
rect 29762 20750 29764 20802
rect 29708 20244 29764 20750
rect 29708 20178 29764 20188
rect 29820 20692 29876 20702
rect 29820 20242 29876 20636
rect 30380 20692 30436 20702
rect 30380 20598 30436 20636
rect 29820 20190 29822 20242
rect 29874 20190 29876 20242
rect 29820 20178 29876 20190
rect 28812 19954 28868 19964
rect 30604 20132 30660 20142
rect 30604 19234 30660 20076
rect 31164 20130 31220 20860
rect 31388 20188 31444 23886
rect 31724 23938 31780 25676
rect 32172 25618 32228 26348
rect 32396 26338 32452 26348
rect 32172 25566 32174 25618
rect 32226 25566 32228 25618
rect 32172 25554 32228 25566
rect 31724 23886 31726 23938
rect 31778 23886 31780 23938
rect 31724 23874 31780 23886
rect 32172 23940 32228 23950
rect 32172 23846 32228 23884
rect 31500 23828 31556 23838
rect 31500 23734 31556 23772
rect 31836 23716 31892 23726
rect 31836 22482 31892 23660
rect 32396 23714 32452 23726
rect 32396 23662 32398 23714
rect 32450 23662 32452 23714
rect 32396 23604 32452 23662
rect 32844 23716 32900 23726
rect 32844 23622 32900 23660
rect 32396 23538 32452 23548
rect 31836 22430 31838 22482
rect 31890 22430 31892 22482
rect 31836 22418 31892 22430
rect 32956 21700 33012 21710
rect 32508 20916 32564 20926
rect 32508 20822 32564 20860
rect 32956 20914 33012 21644
rect 32956 20862 32958 20914
rect 33010 20862 33012 20914
rect 31164 20078 31166 20130
rect 31218 20078 31220 20130
rect 31164 20066 31220 20078
rect 31276 20132 31444 20188
rect 32956 20244 33012 20862
rect 32956 20178 33012 20188
rect 30940 20020 30996 20030
rect 30940 19926 30996 19964
rect 31276 19906 31332 20132
rect 31276 19854 31278 19906
rect 31330 19854 31332 19906
rect 31276 19842 31332 19854
rect 30604 19182 30606 19234
rect 30658 19182 30660 19234
rect 30604 19170 30660 19182
rect 31388 19124 31444 19134
rect 31388 19122 31668 19124
rect 31388 19070 31390 19122
rect 31442 19070 31668 19122
rect 31388 19068 31668 19070
rect 31388 19058 31444 19068
rect 31612 18674 31668 19068
rect 31612 18622 31614 18674
rect 31666 18622 31668 18674
rect 31612 18610 31668 18622
rect 33404 18452 33460 28700
rect 34412 28082 34468 29262
rect 36540 29316 36596 29326
rect 36540 29222 36596 29260
rect 39116 29316 39172 29326
rect 39116 29222 39172 29260
rect 38220 29204 38276 29214
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34972 28756 35028 28766
rect 34972 28662 35028 28700
rect 36316 28420 36372 28430
rect 34412 28030 34414 28082
rect 34466 28030 34468 28082
rect 34412 28018 34468 28030
rect 36092 28418 36372 28420
rect 36092 28366 36318 28418
rect 36370 28366 36372 28418
rect 36092 28364 36372 28366
rect 36092 27970 36148 28364
rect 36316 28354 36372 28364
rect 36092 27918 36094 27970
rect 36146 27918 36148 27970
rect 36092 27906 36148 27918
rect 35308 27860 35364 27870
rect 35084 27858 35364 27860
rect 35084 27806 35310 27858
rect 35362 27806 35364 27858
rect 35084 27804 35364 27806
rect 35084 27076 35140 27804
rect 35308 27794 35364 27804
rect 38220 27746 38276 29148
rect 39228 29204 39284 29214
rect 39228 29110 39284 29148
rect 39788 29202 39844 29214
rect 39788 29150 39790 29202
rect 39842 29150 39844 29202
rect 38892 28420 38948 28430
rect 38220 27694 38222 27746
rect 38274 27694 38276 27746
rect 38220 27682 38276 27694
rect 38668 28418 38948 28420
rect 38668 28366 38894 28418
rect 38946 28366 38948 28418
rect 38668 28364 38948 28366
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 38668 27186 38724 28364
rect 38892 28354 38948 28364
rect 38668 27134 38670 27186
rect 38722 27134 38724 27186
rect 38668 27122 38724 27134
rect 34412 26964 34468 26974
rect 33740 26962 34468 26964
rect 33740 26910 34414 26962
rect 34466 26910 34468 26962
rect 35084 26944 35140 27020
rect 35756 27076 35812 27086
rect 33740 26908 34468 26910
rect 33740 26514 33796 26908
rect 34412 26898 34468 26908
rect 33740 26462 33742 26514
rect 33794 26462 33796 26514
rect 33740 26450 33796 26462
rect 34188 26740 34244 26750
rect 34188 25396 34244 26684
rect 35756 26402 35812 27020
rect 37884 27076 37940 27086
rect 37884 26982 37940 27020
rect 39788 27076 39844 29150
rect 41356 28756 41412 34076
rect 41916 34132 41972 34142
rect 41916 34038 41972 34076
rect 41580 33684 41636 33694
rect 41580 30994 41636 33628
rect 42812 33684 42868 33694
rect 42812 32562 42868 33628
rect 43372 33458 43428 36430
rect 43484 35698 43540 36540
rect 43484 35646 43486 35698
rect 43538 35646 43540 35698
rect 43484 35634 43540 35646
rect 43596 36482 43652 36494
rect 43596 36430 43598 36482
rect 43650 36430 43652 36482
rect 43596 35364 43652 36430
rect 44268 36260 44324 36270
rect 45500 36260 45556 37212
rect 45612 37202 45668 37212
rect 46172 37154 46228 37166
rect 46172 37102 46174 37154
rect 46226 37102 46228 37154
rect 43596 35298 43652 35308
rect 43932 36258 44324 36260
rect 43932 36206 44270 36258
rect 44322 36206 44324 36258
rect 43932 36204 44324 36206
rect 43932 35026 43988 36204
rect 44268 36194 44324 36204
rect 45388 36258 45556 36260
rect 45388 36206 45502 36258
rect 45554 36206 45556 36258
rect 45388 36204 45556 36206
rect 45388 35586 45444 36204
rect 45500 36194 45556 36204
rect 46060 36484 46116 36494
rect 46172 36484 46228 37102
rect 46060 36482 46228 36484
rect 46060 36430 46062 36482
rect 46114 36430 46228 36482
rect 46060 36428 46228 36430
rect 46284 36596 46340 36606
rect 45388 35534 45390 35586
rect 45442 35534 45444 35586
rect 43932 34974 43934 35026
rect 43986 34974 43988 35026
rect 43932 34962 43988 34974
rect 44716 35252 44772 35262
rect 44716 34916 44772 35196
rect 44716 34822 44772 34860
rect 45276 34916 45332 34926
rect 45388 34916 45444 35534
rect 45332 34860 45444 34916
rect 45276 34850 45332 34860
rect 45388 34692 45444 34860
rect 46060 34914 46116 36428
rect 46060 34862 46062 34914
rect 46114 34862 46116 34914
rect 46060 34692 46116 34862
rect 45388 34690 46116 34692
rect 45388 34638 45390 34690
rect 45442 34638 46116 34690
rect 45388 34636 46116 34638
rect 45388 34626 45444 34636
rect 43372 33406 43374 33458
rect 43426 33406 43428 33458
rect 43372 33394 43428 33406
rect 45388 34020 45444 34030
rect 42812 32510 42814 32562
rect 42866 32510 42868 32562
rect 42812 32498 42868 32510
rect 43820 33122 43876 33134
rect 43820 33070 43822 33122
rect 43874 33070 43876 33122
rect 43596 32450 43652 32462
rect 43596 32398 43598 32450
rect 43650 32398 43652 32450
rect 43596 31892 43652 32398
rect 43820 32452 43876 33070
rect 43820 32386 43876 32396
rect 44940 32452 44996 32462
rect 43596 31836 43876 31892
rect 43820 31666 43876 31836
rect 43820 31614 43822 31666
rect 43874 31614 43876 31666
rect 43820 31602 43876 31614
rect 44940 31218 44996 32396
rect 44940 31166 44942 31218
rect 44994 31166 44996 31218
rect 44940 31154 44996 31166
rect 45388 31780 45444 33964
rect 45500 33124 45556 34636
rect 46284 34020 46340 36540
rect 46844 36596 46900 39342
rect 47628 39508 47684 39518
rect 47628 39060 47684 39452
rect 49532 39508 49588 40350
rect 50876 40402 50932 42028
rect 50876 40350 50878 40402
rect 50930 40350 50932 40402
rect 50876 40338 50932 40350
rect 49756 40178 49812 40190
rect 49756 40126 49758 40178
rect 49810 40126 49812 40178
rect 49756 40068 49812 40126
rect 50092 40178 50148 40190
rect 50092 40126 50094 40178
rect 50146 40126 50148 40178
rect 49756 40012 50036 40068
rect 49532 39442 49588 39452
rect 49868 39732 49924 39742
rect 49756 39172 49812 39182
rect 49644 39060 49700 39070
rect 47180 39058 47684 39060
rect 47180 39006 47630 39058
rect 47682 39006 47684 39058
rect 47180 39004 47684 39006
rect 47180 38162 47236 39004
rect 47628 38994 47684 39004
rect 49308 39058 49700 39060
rect 49308 39006 49646 39058
rect 49698 39006 49700 39058
rect 49308 39004 49700 39006
rect 47740 38836 47796 38846
rect 47740 38742 47796 38780
rect 48412 38834 48468 38846
rect 48412 38782 48414 38834
rect 48466 38782 48468 38834
rect 48188 38724 48244 38734
rect 47180 38110 47182 38162
rect 47234 38110 47236 38162
rect 47180 38098 47236 38110
rect 47852 38610 47908 38622
rect 47852 38558 47854 38610
rect 47906 38558 47908 38610
rect 47852 37156 47908 38558
rect 48188 38500 48244 38668
rect 48188 37266 48244 38444
rect 48188 37214 48190 37266
rect 48242 37214 48244 37266
rect 48188 37202 48244 37214
rect 48412 37268 48468 38782
rect 48412 37202 48468 37212
rect 48524 38722 48580 38734
rect 48524 38670 48526 38722
rect 48578 38670 48580 38722
rect 48524 37266 48580 38670
rect 48748 38612 48804 38622
rect 48748 38518 48804 38556
rect 49308 38162 49364 39004
rect 49644 38994 49700 39004
rect 49532 38836 49588 38846
rect 49532 38742 49588 38780
rect 49756 38834 49812 39116
rect 49756 38782 49758 38834
rect 49810 38782 49812 38834
rect 49756 38770 49812 38782
rect 49308 38110 49310 38162
rect 49362 38110 49364 38162
rect 49308 38098 49364 38110
rect 49756 38612 49812 38622
rect 48524 37214 48526 37266
rect 48578 37214 48580 37266
rect 48524 37202 48580 37214
rect 48972 37268 49028 37278
rect 47852 37090 47908 37100
rect 46844 36530 46900 36540
rect 46956 37044 47012 37054
rect 46844 36372 46900 36382
rect 46956 36372 47012 36988
rect 48076 37044 48132 37054
rect 48076 36950 48132 36988
rect 48412 37044 48468 37054
rect 48412 36950 48468 36988
rect 48972 36594 49028 37212
rect 49532 37268 49588 37278
rect 49532 37174 49588 37212
rect 49756 37268 49812 38556
rect 49756 37136 49812 37212
rect 49868 38052 49924 39676
rect 49980 38836 50036 40012
rect 50092 39172 50148 40126
rect 51212 39620 51268 43372
rect 52332 42868 52388 43596
rect 53004 43652 53060 45052
rect 54012 44324 54068 44334
rect 54124 44324 54180 46510
rect 54460 44324 54516 44334
rect 54124 44322 54516 44324
rect 54124 44270 54462 44322
rect 54514 44270 54516 44322
rect 54124 44268 54516 44270
rect 54012 44230 54068 44268
rect 54460 44258 54516 44268
rect 53452 44212 53508 44222
rect 53004 43586 53060 43596
rect 53228 44210 53508 44212
rect 53228 44158 53454 44210
rect 53506 44158 53508 44210
rect 53228 44156 53508 44158
rect 53228 43204 53284 44156
rect 53452 44146 53508 44156
rect 51884 42866 52388 42868
rect 51884 42814 52334 42866
rect 52386 42814 52388 42866
rect 51884 42812 52388 42814
rect 51884 42756 51940 42812
rect 52332 42802 52388 42812
rect 52892 43148 53284 43204
rect 53340 43652 53396 43662
rect 51884 42624 51940 42700
rect 52892 41858 52948 43148
rect 53340 42196 53396 43596
rect 53340 42064 53396 42140
rect 54124 42196 54180 42206
rect 52892 41806 52894 41858
rect 52946 41806 52948 41858
rect 52892 41794 52948 41806
rect 54124 40626 54180 42140
rect 54124 40574 54126 40626
rect 54178 40574 54180 40626
rect 54124 40562 54180 40574
rect 51548 40292 51604 40302
rect 51212 39526 51268 39564
rect 51324 40290 51604 40292
rect 51324 40238 51550 40290
rect 51602 40238 51604 40290
rect 51324 40236 51604 40238
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50092 39106 50148 39116
rect 51212 39060 51268 39070
rect 49980 38780 50148 38836
rect 49980 38610 50036 38622
rect 49980 38558 49982 38610
rect 50034 38558 50036 38610
rect 49980 38500 50036 38558
rect 49980 38434 50036 38444
rect 49980 38052 50036 38062
rect 49868 38050 50036 38052
rect 49868 37998 49982 38050
rect 50034 37998 50036 38050
rect 49868 37996 50036 37998
rect 48972 36542 48974 36594
rect 49026 36542 49028 36594
rect 48972 36530 49028 36542
rect 49868 36482 49924 37996
rect 49980 37986 50036 37996
rect 50092 37490 50148 38780
rect 51212 38834 51268 39004
rect 51324 39058 51380 40236
rect 51548 40226 51604 40236
rect 53676 40292 53732 40302
rect 53676 40290 54068 40292
rect 53676 40238 53678 40290
rect 53730 40238 54068 40290
rect 53676 40236 54068 40238
rect 53676 40226 53732 40236
rect 53676 39732 53732 39742
rect 53676 39638 53732 39676
rect 51324 39006 51326 39058
rect 51378 39006 51380 39058
rect 51324 38994 51380 39006
rect 52332 39620 52388 39630
rect 52332 39058 52388 39564
rect 53452 39508 53508 39518
rect 52332 39006 52334 39058
rect 52386 39006 52388 39058
rect 52332 38948 52388 39006
rect 52332 38882 52388 38892
rect 53004 39506 53508 39508
rect 53004 39454 53454 39506
rect 53506 39454 53508 39506
rect 53004 39452 53508 39454
rect 51212 38782 51214 38834
rect 51266 38782 51268 38834
rect 51212 38770 51268 38782
rect 51660 38836 51716 38846
rect 51660 38742 51716 38780
rect 52444 38836 52500 38846
rect 50988 38724 51044 38734
rect 50652 38500 50708 38510
rect 50652 38050 50708 38444
rect 50652 37998 50654 38050
rect 50706 37998 50708 38050
rect 50652 37986 50708 37998
rect 50988 37938 51044 38668
rect 51436 38724 51492 38734
rect 52444 38668 52500 38780
rect 51436 38630 51492 38668
rect 52332 38612 52500 38668
rect 53004 38834 53060 39452
rect 53452 39442 53508 39452
rect 53676 39508 53732 39518
rect 53676 39414 53732 39452
rect 53004 38782 53006 38834
rect 53058 38782 53060 38834
rect 53004 38724 53060 38782
rect 53452 38948 53508 38958
rect 53004 38658 53060 38668
rect 53340 38724 53396 38734
rect 53340 38630 53396 38668
rect 52892 38612 52948 38622
rect 52108 38164 52164 38174
rect 52108 38070 52164 38108
rect 50988 37886 50990 37938
rect 51042 37886 51044 37938
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50092 37438 50094 37490
rect 50146 37438 50148 37490
rect 50092 37044 50148 37438
rect 50988 37268 51044 37886
rect 52332 38050 52388 38612
rect 52892 38518 52948 38556
rect 53228 38610 53284 38622
rect 53228 38558 53230 38610
rect 53282 38558 53284 38610
rect 53228 38388 53284 38558
rect 52668 38332 53284 38388
rect 52668 38274 52724 38332
rect 52668 38222 52670 38274
rect 52722 38222 52724 38274
rect 52668 38210 52724 38222
rect 52332 37998 52334 38050
rect 52386 37998 52388 38050
rect 52332 37604 52388 37998
rect 52780 38164 52836 38174
rect 52332 37548 52724 37604
rect 52556 37380 52612 37390
rect 51100 37268 51156 37278
rect 50988 37266 51156 37268
rect 50988 37214 51102 37266
rect 51154 37214 51156 37266
rect 50988 37212 51156 37214
rect 51100 37202 51156 37212
rect 51324 37268 51380 37278
rect 51324 37174 51380 37212
rect 51548 37268 51604 37278
rect 51548 37174 51604 37212
rect 52108 37156 52164 37166
rect 52108 37062 52164 37100
rect 50988 37044 51044 37054
rect 50092 36978 50148 36988
rect 50540 37042 51044 37044
rect 50540 36990 50990 37042
rect 51042 36990 51044 37042
rect 50540 36988 51044 36990
rect 50540 36594 50596 36988
rect 50988 36978 51044 36988
rect 50540 36542 50542 36594
rect 50594 36542 50596 36594
rect 50540 36530 50596 36542
rect 52556 36596 52612 37324
rect 52668 37378 52724 37548
rect 52668 37326 52670 37378
rect 52722 37326 52724 37378
rect 52668 37314 52724 37326
rect 52780 37378 52836 38108
rect 52780 37326 52782 37378
rect 52834 37326 52836 37378
rect 52780 37314 52836 37326
rect 53228 37380 53284 38332
rect 53452 38050 53508 38892
rect 54012 38946 54068 40236
rect 54572 39732 54628 46620
rect 54684 46564 54740 46574
rect 54684 44434 54740 46508
rect 54684 44382 54686 44434
rect 54738 44382 54740 44434
rect 54684 44370 54740 44382
rect 55132 44996 55188 45006
rect 55132 44210 55188 44940
rect 55916 44996 55972 45006
rect 55916 44902 55972 44940
rect 56364 44994 56420 45006
rect 56364 44942 56366 44994
rect 56418 44942 56420 44994
rect 55132 44158 55134 44210
rect 55186 44158 55188 44210
rect 55132 44146 55188 44158
rect 56364 43708 56420 44942
rect 56252 43652 56420 43708
rect 56252 43520 56308 43596
rect 54572 39666 54628 39676
rect 54012 38894 54014 38946
rect 54066 38894 54068 38946
rect 54012 38836 54068 38894
rect 54012 38770 54068 38780
rect 54348 38834 54404 38846
rect 54348 38782 54350 38834
rect 54402 38782 54404 38834
rect 54124 38724 54180 38734
rect 54124 38630 54180 38668
rect 54236 38612 54292 38622
rect 54236 38162 54292 38556
rect 54236 38110 54238 38162
rect 54290 38110 54292 38162
rect 54236 38098 54292 38110
rect 54348 38164 54404 38782
rect 54348 38098 54404 38108
rect 56364 38164 56420 38174
rect 56364 38070 56420 38108
rect 53452 37998 53454 38050
rect 53506 37998 53508 38050
rect 53452 37986 53508 37998
rect 53452 37380 53508 37390
rect 53228 37378 53508 37380
rect 53228 37326 53454 37378
rect 53506 37326 53508 37378
rect 53228 37324 53508 37326
rect 53452 37314 53508 37324
rect 53676 37380 53732 37390
rect 53676 37286 53732 37324
rect 53564 37268 53620 37278
rect 53564 37174 53620 37212
rect 52668 36596 52724 36606
rect 52556 36594 52724 36596
rect 52556 36542 52670 36594
rect 52722 36542 52724 36594
rect 52556 36540 52724 36542
rect 52668 36530 52724 36540
rect 49868 36430 49870 36482
rect 49922 36430 49924 36482
rect 49868 36418 49924 36430
rect 46844 36370 47012 36372
rect 46844 36318 46846 36370
rect 46898 36318 47012 36370
rect 46844 36316 47012 36318
rect 46844 36306 46900 36316
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 48076 35586 48132 35598
rect 48076 35534 48078 35586
rect 48130 35534 48132 35586
rect 46844 34802 46900 34814
rect 46844 34750 46846 34802
rect 46898 34750 46900 34802
rect 46844 34356 46900 34750
rect 46844 34290 46900 34300
rect 47740 34356 47796 34366
rect 47740 34262 47796 34300
rect 46284 33954 46340 33964
rect 48076 34020 48132 35534
rect 48076 33954 48132 33964
rect 48972 35026 49028 35038
rect 48972 34974 48974 35026
rect 49026 34974 49028 35026
rect 45724 33124 45780 33134
rect 45500 33122 45780 33124
rect 45500 33070 45726 33122
rect 45778 33070 45780 33122
rect 45500 33068 45780 33070
rect 45612 32452 45668 33068
rect 45724 33058 45780 33068
rect 46844 32674 46900 32686
rect 46844 32622 46846 32674
rect 46898 32622 46900 32674
rect 45612 32386 45668 32396
rect 45724 32450 45780 32462
rect 45724 32398 45726 32450
rect 45778 32398 45780 32450
rect 45724 31948 45780 32398
rect 46172 32452 46228 32462
rect 46172 32358 46228 32396
rect 46844 31948 46900 32622
rect 41580 30942 41582 30994
rect 41634 30942 41636 30994
rect 41580 30930 41636 30942
rect 42364 30884 42420 30894
rect 44492 30884 44548 30894
rect 42364 30882 43540 30884
rect 42364 30830 42366 30882
rect 42418 30830 43540 30882
rect 42364 30828 43540 30830
rect 42364 30818 42420 30828
rect 43484 30098 43540 30828
rect 44492 30882 45220 30884
rect 44492 30830 44494 30882
rect 44546 30830 45220 30882
rect 44492 30828 45220 30830
rect 44492 30818 44548 30828
rect 44156 30212 44212 30222
rect 44156 30118 44212 30156
rect 43484 30046 43486 30098
rect 43538 30046 43540 30098
rect 43484 30034 43540 30046
rect 41580 29428 41636 29438
rect 41580 29334 41636 29372
rect 45164 29426 45220 30828
rect 45388 30212 45444 31724
rect 45388 30146 45444 30156
rect 45612 31892 45780 31948
rect 46620 31892 46900 31948
rect 48972 31948 49028 34974
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 49868 32674 49924 32686
rect 49868 32622 49870 32674
rect 49922 32622 49924 32674
rect 49868 31948 49924 32622
rect 48972 31892 49364 31948
rect 49868 31892 50372 31948
rect 45164 29374 45166 29426
rect 45218 29374 45220 29426
rect 45164 29362 45220 29374
rect 45612 29426 45668 31892
rect 46620 31106 46676 31892
rect 46844 31780 46900 31790
rect 46844 31686 46900 31724
rect 46620 31054 46622 31106
rect 46674 31054 46676 31106
rect 46620 31042 46676 31054
rect 45948 30996 46004 31006
rect 45724 30940 45948 30996
rect 45724 30210 45780 30940
rect 45948 30902 46004 30940
rect 48748 30884 48804 30894
rect 48748 30882 49140 30884
rect 48748 30830 48750 30882
rect 48802 30830 49140 30882
rect 48748 30828 49140 30830
rect 48748 30818 48804 30828
rect 48524 30324 48580 30334
rect 48524 30230 48580 30268
rect 45724 30158 45726 30210
rect 45778 30158 45780 30210
rect 45724 30146 45780 30158
rect 49084 30210 49140 30828
rect 49308 30434 49364 31892
rect 49532 31666 49588 31678
rect 49532 31614 49534 31666
rect 49586 31614 49588 31666
rect 49532 30996 49588 31614
rect 50316 31106 50372 31892
rect 51212 31780 51268 31790
rect 51212 31686 51268 31724
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50316 31054 50318 31106
rect 50370 31054 50372 31106
rect 50316 31042 50372 31054
rect 49532 30864 49588 30940
rect 52444 30882 52500 30894
rect 52444 30830 52446 30882
rect 52498 30830 52500 30882
rect 49308 30382 49310 30434
rect 49362 30382 49364 30434
rect 49308 30370 49364 30382
rect 49756 30436 49812 30446
rect 49756 30342 49812 30380
rect 52444 30436 52500 30830
rect 52444 30370 52500 30380
rect 49532 30324 49588 30334
rect 49532 30230 49588 30268
rect 49084 30158 49086 30210
rect 49138 30158 49140 30210
rect 49084 30146 49140 30158
rect 46396 30098 46452 30110
rect 46396 30046 46398 30098
rect 46450 30046 46452 30098
rect 46396 29652 46452 30046
rect 49644 29986 49700 29998
rect 49644 29934 49646 29986
rect 49698 29934 49700 29986
rect 46508 29652 46564 29662
rect 46396 29650 46564 29652
rect 46396 29598 46510 29650
rect 46562 29598 46564 29650
rect 46396 29596 46564 29598
rect 46508 29586 46564 29596
rect 45612 29374 45614 29426
rect 45666 29374 45668 29426
rect 45612 29362 45668 29374
rect 49644 29428 49700 29934
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 49756 29428 49812 29438
rect 49644 29426 49812 29428
rect 49644 29374 49758 29426
rect 49810 29374 49812 29426
rect 49644 29372 49812 29374
rect 49756 29362 49812 29372
rect 41356 28690 41412 28700
rect 42364 29314 42420 29326
rect 42364 29262 42366 29314
rect 42418 29262 42420 29314
rect 42252 28532 42308 28542
rect 42364 28532 42420 29262
rect 44492 29316 44548 29326
rect 44492 29222 44548 29260
rect 45388 29316 45444 29326
rect 45388 29222 45444 29260
rect 45948 29316 46004 29326
rect 45948 29222 46004 29260
rect 49532 29316 49588 29326
rect 49532 29222 49588 29260
rect 42252 28530 42420 28532
rect 42252 28478 42254 28530
rect 42306 28478 42420 28530
rect 42252 28476 42420 28478
rect 45836 29202 45892 29214
rect 45836 29150 45838 29202
rect 45890 29150 45892 29202
rect 45836 28532 45892 29150
rect 50092 29202 50148 29214
rect 50092 29150 50094 29202
rect 50146 29150 50148 29202
rect 49756 28642 49812 28654
rect 49756 28590 49758 28642
rect 49810 28590 49812 28642
rect 45836 28476 46340 28532
rect 42252 28466 42308 28476
rect 44268 28418 44324 28430
rect 44268 28366 44270 28418
rect 44322 28366 44324 28418
rect 41580 27972 41636 27982
rect 40908 27970 41636 27972
rect 40908 27918 41582 27970
rect 41634 27918 41636 27970
rect 40908 27916 41636 27918
rect 39788 27010 39844 27020
rect 40796 27186 40852 27198
rect 40796 27134 40798 27186
rect 40850 27134 40852 27186
rect 35756 26350 35758 26402
rect 35810 26350 35812 26402
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 34300 25620 34356 25630
rect 34300 25618 34692 25620
rect 34300 25566 34302 25618
rect 34354 25566 34692 25618
rect 34300 25564 34692 25566
rect 34300 25554 34356 25564
rect 34188 25340 34468 25396
rect 34412 24162 34468 25340
rect 34412 24110 34414 24162
rect 34466 24110 34468 24162
rect 34412 24098 34468 24110
rect 34636 24162 34692 25564
rect 34636 24110 34638 24162
rect 34690 24110 34692 24162
rect 34636 24098 34692 24110
rect 34748 25508 34804 25518
rect 34300 23940 34356 23950
rect 34300 23846 34356 23884
rect 33628 23044 33684 23054
rect 33628 22950 33684 22988
rect 33964 22708 34020 22718
rect 33964 22482 34020 22652
rect 33964 22430 33966 22482
rect 34018 22430 34020 22482
rect 33964 22418 34020 22430
rect 34748 22484 34804 25452
rect 35756 24724 35812 26350
rect 40236 26292 40292 26302
rect 40236 26198 40292 26236
rect 40796 26180 40852 27134
rect 40796 26114 40852 26124
rect 39788 26068 39844 26078
rect 38108 25452 38388 25508
rect 37660 25396 37716 25406
rect 38108 25396 38164 25452
rect 37660 25394 38164 25396
rect 37660 25342 37662 25394
rect 37714 25342 38164 25394
rect 37660 25340 38164 25342
rect 37660 25330 37716 25340
rect 38220 25284 38276 25294
rect 37772 25282 38276 25284
rect 37772 25230 38222 25282
rect 38274 25230 38276 25282
rect 37772 25228 38276 25230
rect 37772 24948 37828 25228
rect 38220 25218 38276 25228
rect 36988 24892 37828 24948
rect 36988 24834 37044 24892
rect 36988 24782 36990 24834
rect 37042 24782 37044 24834
rect 36988 24770 37044 24782
rect 36204 24724 36260 24734
rect 35756 24722 36260 24724
rect 35756 24670 36206 24722
rect 36258 24670 36260 24722
rect 35756 24668 36260 24670
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34860 23938 34916 23950
rect 34860 23886 34862 23938
rect 34914 23886 34916 23938
rect 34860 23044 34916 23886
rect 34860 22978 34916 22988
rect 34972 23938 35028 23950
rect 34972 23886 34974 23938
rect 35026 23886 35028 23938
rect 34972 22708 35028 23886
rect 36204 23940 36260 24668
rect 38332 24050 38388 25452
rect 39676 24836 39732 24846
rect 38332 23998 38334 24050
rect 38386 23998 38388 24050
rect 38332 23986 38388 23998
rect 38780 24834 39732 24836
rect 38780 24782 39678 24834
rect 39730 24782 39732 24834
rect 38780 24780 39732 24782
rect 36204 23874 36260 23884
rect 36540 23940 36596 23950
rect 36540 23154 36596 23884
rect 37548 23940 37604 23950
rect 37548 23846 37604 23884
rect 38668 23716 38724 23726
rect 36540 23102 36542 23154
rect 36594 23102 36596 23154
rect 36540 23090 36596 23102
rect 36764 23604 36820 23614
rect 35756 23042 35812 23054
rect 35756 22990 35758 23042
rect 35810 22990 35812 23042
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 34972 22642 35028 22652
rect 35084 22484 35140 22494
rect 34748 22482 35140 22484
rect 34748 22430 35086 22482
rect 35138 22430 35140 22482
rect 34748 22428 35140 22430
rect 34636 22260 34692 22270
rect 34636 22166 34692 22204
rect 33740 21700 33796 21710
rect 33740 20802 33796 21644
rect 35084 21700 35140 22428
rect 35756 22260 35812 22990
rect 35756 22194 35812 22204
rect 35084 21634 35140 21644
rect 35644 21700 35700 21710
rect 35644 21606 35700 21644
rect 34972 21588 35028 21598
rect 34972 21494 35028 21532
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 33740 20750 33742 20802
rect 33794 20750 33796 20802
rect 33740 20188 33796 20750
rect 36540 20914 36596 20926
rect 36540 20862 36542 20914
rect 36594 20862 36596 20914
rect 34412 20690 34468 20702
rect 34412 20638 34414 20690
rect 34466 20638 34468 20690
rect 33964 20244 34020 20254
rect 33740 20132 34020 20188
rect 34300 20244 34356 20254
rect 34412 20244 34468 20638
rect 35644 20580 35700 20590
rect 34300 20242 34468 20244
rect 34300 20190 34302 20242
rect 34354 20190 34468 20242
rect 34300 20188 34468 20190
rect 34860 20244 34916 20254
rect 34300 20178 34356 20188
rect 33404 18386 33460 18396
rect 33516 19346 33572 19358
rect 33516 19294 33518 19346
rect 33570 19294 33572 19346
rect 28588 18338 28644 18350
rect 28588 18286 28590 18338
rect 28642 18286 28644 18338
rect 27580 17108 27636 17118
rect 27580 17014 27636 17052
rect 28140 17108 28196 17118
rect 28140 16882 28196 17052
rect 28140 16830 28142 16882
rect 28194 16830 28196 16882
rect 28140 16818 28196 16830
rect 27132 15876 27188 15886
rect 26908 15874 27188 15876
rect 26908 15822 27134 15874
rect 27186 15822 27188 15874
rect 26908 15820 27188 15822
rect 26908 15426 26964 15820
rect 27132 15810 27188 15820
rect 26908 15374 26910 15426
rect 26962 15374 26964 15426
rect 26908 15362 26964 15374
rect 26796 14924 26964 14980
rect 26908 13746 26964 14924
rect 26908 13694 26910 13746
rect 26962 13694 26964 13746
rect 26908 13682 26964 13694
rect 27916 14644 27972 14654
rect 26236 13458 26292 13468
rect 27916 13186 27972 14588
rect 28140 14642 28196 14654
rect 28140 14590 28142 14642
rect 28194 14590 28196 14642
rect 27916 13134 27918 13186
rect 27970 13134 27972 13186
rect 27916 13122 27972 13134
rect 28028 13188 28084 13198
rect 28140 13188 28196 14590
rect 28588 13412 28644 18286
rect 29036 18338 29092 18350
rect 29036 18286 29038 18338
rect 29090 18286 29092 18338
rect 29036 17108 29092 18286
rect 33516 18340 33572 19294
rect 33852 19012 33908 20132
rect 34860 20018 34916 20188
rect 35644 20130 35700 20524
rect 35644 20078 35646 20130
rect 35698 20078 35700 20130
rect 35644 20066 35700 20078
rect 36540 20132 36596 20862
rect 36540 20066 36596 20076
rect 34860 19966 34862 20018
rect 34914 19966 34916 20018
rect 34860 19954 34916 19966
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 33964 19012 34020 19022
rect 33852 19010 34132 19012
rect 33852 18958 33966 19010
rect 34018 18958 34132 19010
rect 33852 18956 34132 18958
rect 33964 18946 34020 18956
rect 34076 18450 34132 18956
rect 34076 18398 34078 18450
rect 34130 18398 34132 18450
rect 34076 18386 34132 18398
rect 33516 18274 33572 18284
rect 34636 18340 34692 18350
rect 29596 17444 29652 17454
rect 29036 17042 29092 17052
rect 29148 17442 29652 17444
rect 29148 17390 29598 17442
rect 29650 17390 29652 17442
rect 29148 17388 29652 17390
rect 28924 16884 28980 16894
rect 29148 16884 29204 17388
rect 29596 17378 29652 17388
rect 31612 16996 31668 17006
rect 31164 16994 31668 16996
rect 31164 16942 31614 16994
rect 31666 16942 31668 16994
rect 31164 16940 31668 16942
rect 28924 16882 29204 16884
rect 28924 16830 28926 16882
rect 28978 16830 29204 16882
rect 28924 16828 29204 16830
rect 31052 16884 31108 16894
rect 28924 16818 28980 16828
rect 31052 16770 31108 16828
rect 31052 16718 31054 16770
rect 31106 16718 31108 16770
rect 31052 16706 31108 16718
rect 31164 16436 31220 16940
rect 31612 16930 31668 16940
rect 32956 16996 33012 17006
rect 30828 16380 31220 16436
rect 30828 16210 30884 16380
rect 30828 16158 30830 16210
rect 30882 16158 30884 16210
rect 30828 16146 30884 16158
rect 32956 16210 33012 16940
rect 33740 16996 33796 17006
rect 33740 16902 33796 16940
rect 33628 16884 33684 16894
rect 33628 16790 33684 16828
rect 34636 16882 34692 18284
rect 34860 18340 34916 18350
rect 34860 18338 35140 18340
rect 34860 18286 34862 18338
rect 34914 18286 35140 18338
rect 34860 18284 35140 18286
rect 34860 18274 34916 18284
rect 35084 17554 35140 18284
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35084 17502 35086 17554
rect 35138 17502 35140 17554
rect 35084 17490 35140 17502
rect 34748 17108 34804 17118
rect 34748 17014 34804 17052
rect 36764 17106 36820 23548
rect 38668 23266 38724 23660
rect 38668 23214 38670 23266
rect 38722 23214 38724 23266
rect 38668 23202 38724 23214
rect 37996 23154 38052 23166
rect 37996 23102 37998 23154
rect 38050 23102 38052 23154
rect 37996 22372 38052 23102
rect 38668 22484 38724 22494
rect 38780 22484 38836 24780
rect 39676 24770 39732 24780
rect 39116 24612 39172 24622
rect 39788 24612 39844 26012
rect 40796 25620 40852 25630
rect 40908 25620 40964 27916
rect 41580 27906 41636 27916
rect 44156 27972 44212 27982
rect 44268 27972 44324 28366
rect 44156 27970 44324 27972
rect 44156 27918 44158 27970
rect 44210 27918 44324 27970
rect 44156 27916 44324 27918
rect 44156 27906 44212 27916
rect 43484 27860 43540 27870
rect 43484 27766 43540 27804
rect 46284 27746 46340 28476
rect 49308 28418 49364 28430
rect 49308 28366 49310 28418
rect 49362 28366 49364 28418
rect 46284 27694 46286 27746
rect 46338 27694 46340 27746
rect 46284 27682 46340 27694
rect 46508 27860 46564 27870
rect 41804 27076 41860 27086
rect 41804 26982 41860 27020
rect 46508 27074 46564 27804
rect 46732 27860 46788 27870
rect 46732 27766 46788 27804
rect 48076 27860 48132 27870
rect 49308 27860 49364 28366
rect 49532 27860 49588 27870
rect 49308 27858 49588 27860
rect 49308 27806 49534 27858
rect 49586 27806 49588 27858
rect 49308 27804 49588 27806
rect 48076 27766 48132 27804
rect 48748 27748 48804 27758
rect 48748 27746 49252 27748
rect 48748 27694 48750 27746
rect 48802 27694 49252 27746
rect 48748 27692 49252 27694
rect 48748 27682 48804 27692
rect 48636 27636 48692 27646
rect 46508 27022 46510 27074
rect 46562 27022 46564 27074
rect 46508 27010 46564 27022
rect 48524 27634 48692 27636
rect 48524 27582 48638 27634
rect 48690 27582 48692 27634
rect 48524 27580 48692 27582
rect 41692 26962 41748 26974
rect 41692 26910 41694 26962
rect 41746 26910 41748 26962
rect 41580 26292 41636 26302
rect 40796 25618 40964 25620
rect 40796 25566 40798 25618
rect 40850 25566 40964 25618
rect 40796 25564 40964 25566
rect 41020 26290 41636 26292
rect 41020 26238 41582 26290
rect 41634 26238 41636 26290
rect 41020 26236 41636 26238
rect 40796 25554 40852 25564
rect 40124 25508 40180 25518
rect 40124 25414 40180 25452
rect 39116 24610 39844 24612
rect 39116 24558 39118 24610
rect 39170 24558 39844 24610
rect 39116 24556 39844 24558
rect 39116 24546 39172 24556
rect 41020 24500 41076 26236
rect 41580 26226 41636 26236
rect 40460 24444 41076 24500
rect 40460 24050 40516 24444
rect 40460 23998 40462 24050
rect 40514 23998 40516 24050
rect 40460 23986 40516 23998
rect 41020 23716 41076 23726
rect 41020 23622 41076 23660
rect 40796 23044 40852 23054
rect 38668 22482 38836 22484
rect 38668 22430 38670 22482
rect 38722 22430 38836 22482
rect 38668 22428 38836 22430
rect 40684 23042 40852 23044
rect 40684 22990 40798 23042
rect 40850 22990 40852 23042
rect 40684 22988 40852 22990
rect 38668 22418 38724 22428
rect 37996 22240 38052 22316
rect 39228 22372 39284 22382
rect 39228 21700 39284 22316
rect 40684 22260 40740 22988
rect 40796 22978 40852 22988
rect 41580 22596 41636 22606
rect 40796 22594 41636 22596
rect 40796 22542 41582 22594
rect 41634 22542 41636 22594
rect 40796 22540 41636 22542
rect 41692 22596 41748 26910
rect 41916 26962 41972 26974
rect 41916 26910 41918 26962
rect 41970 26910 41972 26962
rect 41916 26516 41972 26910
rect 47180 26964 47236 26974
rect 48524 26964 48580 27580
rect 48636 27570 48692 27580
rect 49196 27188 49252 27692
rect 49308 27188 49364 27198
rect 49196 27186 49364 27188
rect 49196 27134 49310 27186
rect 49362 27134 49364 27186
rect 49196 27132 49364 27134
rect 49308 27122 49364 27132
rect 47180 26962 48468 26964
rect 47180 26910 47182 26962
rect 47234 26910 48468 26962
rect 47180 26908 48468 26910
rect 47180 26898 47236 26908
rect 42364 26850 42420 26862
rect 42364 26798 42366 26850
rect 42418 26798 42420 26850
rect 42140 26516 42196 26526
rect 41916 26514 42196 26516
rect 41916 26462 42142 26514
rect 42194 26462 42196 26514
rect 41916 26460 42196 26462
rect 42140 26450 42196 26460
rect 42364 26516 42420 26798
rect 42364 26450 42420 26460
rect 48412 26514 48468 26908
rect 48412 26462 48414 26514
rect 48466 26462 48468 26514
rect 48412 26450 48468 26462
rect 42252 26292 42308 26302
rect 42812 26292 42868 26302
rect 42252 26290 42644 26292
rect 42252 26238 42254 26290
rect 42306 26238 42644 26290
rect 42252 26236 42644 26238
rect 42252 26226 42308 26236
rect 42028 26180 42084 26190
rect 42028 26086 42084 26124
rect 41804 26068 41860 26078
rect 41804 25974 41860 26012
rect 42588 26066 42644 26236
rect 42588 26014 42590 26066
rect 42642 26014 42644 26066
rect 42588 26002 42644 26014
rect 42812 26178 42868 26236
rect 43596 26292 43652 26302
rect 43596 26290 43764 26292
rect 43596 26238 43598 26290
rect 43650 26238 43764 26290
rect 43596 26236 43764 26238
rect 43596 26226 43652 26236
rect 42812 26126 42814 26178
rect 42866 26126 42868 26178
rect 41804 25508 41860 25518
rect 41804 24836 41860 25452
rect 41804 23938 41860 24780
rect 42588 24612 42644 24622
rect 42588 24050 42644 24556
rect 42588 23998 42590 24050
rect 42642 23998 42644 24050
rect 42588 23986 42644 23998
rect 41804 23886 41806 23938
rect 41858 23886 41860 23938
rect 41804 23874 41860 23886
rect 42028 23156 42084 23166
rect 41916 22596 41972 22606
rect 41692 22594 41972 22596
rect 41692 22542 41918 22594
rect 41970 22542 41972 22594
rect 41692 22540 41972 22542
rect 40796 22482 40852 22540
rect 41580 22530 41636 22540
rect 41916 22530 41972 22540
rect 40796 22430 40798 22482
rect 40850 22430 40852 22482
rect 40796 22418 40852 22430
rect 41356 22370 41412 22382
rect 41356 22318 41358 22370
rect 41410 22318 41412 22370
rect 41356 22260 41412 22318
rect 41804 22372 41860 22382
rect 41804 22370 41972 22372
rect 41804 22318 41806 22370
rect 41858 22318 41972 22370
rect 41804 22316 41972 22318
rect 41804 22306 41860 22316
rect 40684 22204 41412 22260
rect 39228 20802 39284 21644
rect 41468 21700 41524 21710
rect 39340 21588 39396 21598
rect 39340 21494 39396 21532
rect 39228 20750 39230 20802
rect 39282 20750 39284 20802
rect 39228 20738 39284 20750
rect 40012 20690 40068 20702
rect 40012 20638 40014 20690
rect 40066 20638 40068 20690
rect 37548 20580 37604 20590
rect 37548 20486 37604 20524
rect 38108 20580 38164 20590
rect 38556 20580 38612 20590
rect 38108 20578 38612 20580
rect 38108 20526 38110 20578
rect 38162 20526 38558 20578
rect 38610 20526 38612 20578
rect 38108 20524 38612 20526
rect 37436 20244 37492 20254
rect 36988 20020 37044 20030
rect 36988 18338 37044 19964
rect 37436 18450 37492 20188
rect 38108 20244 38164 20524
rect 38556 20514 38612 20524
rect 38108 20178 38164 20188
rect 38556 20242 38612 20254
rect 38556 20190 38558 20242
rect 38610 20190 38612 20242
rect 38444 20132 38500 20142
rect 38444 20038 38500 20076
rect 38332 20020 38388 20030
rect 38332 19926 38388 19964
rect 37772 19908 37828 19918
rect 37772 19814 37828 19852
rect 38108 19236 38164 19246
rect 38108 19142 38164 19180
rect 38556 18564 38612 20190
rect 40012 20244 40068 20638
rect 40012 20178 40068 20188
rect 40572 20244 40628 20282
rect 40572 20178 40628 20188
rect 39900 20130 39956 20142
rect 39900 20078 39902 20130
rect 39954 20078 39956 20130
rect 39340 20018 39396 20030
rect 39340 19966 39342 20018
rect 39394 19966 39396 20018
rect 39340 19908 39396 19966
rect 39340 19842 39396 19852
rect 39900 19348 39956 20078
rect 41468 20132 41524 21644
rect 41916 21364 41972 22316
rect 42028 21588 42084 23100
rect 42812 23156 42868 26126
rect 42924 26066 42980 26078
rect 42924 26014 42926 26066
rect 42978 26014 42980 26066
rect 42924 25618 42980 26014
rect 42924 25566 42926 25618
rect 42978 25566 42980 25618
rect 42924 25554 42980 25566
rect 43372 25284 43428 25294
rect 43708 25284 43764 26236
rect 48076 26290 48132 26302
rect 48076 26238 48078 26290
rect 48130 26238 48132 26290
rect 44268 26178 44324 26190
rect 46396 26180 46452 26190
rect 44268 26126 44270 26178
rect 44322 26126 44324 26178
rect 44268 25732 44324 26126
rect 45948 26178 46452 26180
rect 45948 26126 46398 26178
rect 46450 26126 46452 26178
rect 45948 26124 46452 26126
rect 45948 25844 46004 26124
rect 46396 26114 46452 26124
rect 46844 26178 46900 26190
rect 46844 26126 46846 26178
rect 46898 26126 46900 26178
rect 45724 25788 46004 25844
rect 44380 25732 44436 25742
rect 44268 25730 44436 25732
rect 44268 25678 44382 25730
rect 44434 25678 44436 25730
rect 44268 25676 44436 25678
rect 44380 25666 44436 25676
rect 44716 25396 44772 25406
rect 44716 25302 44772 25340
rect 45500 25396 45556 25406
rect 45500 25302 45556 25340
rect 43372 25282 43764 25284
rect 43372 25230 43374 25282
rect 43426 25230 43764 25282
rect 43372 25228 43764 25230
rect 43372 25218 43428 25228
rect 43708 24948 43764 25228
rect 44492 25284 44548 25294
rect 44492 25190 44548 25228
rect 45388 25284 45444 25294
rect 43708 24882 43764 24892
rect 44940 24948 44996 24958
rect 44716 24052 44772 24062
rect 44716 23958 44772 23996
rect 44940 23268 44996 24892
rect 45388 24836 45444 25228
rect 45500 24836 45556 24846
rect 45388 24834 45556 24836
rect 45388 24782 45502 24834
rect 45554 24782 45556 24834
rect 45388 24780 45556 24782
rect 45500 24770 45556 24780
rect 45612 24612 45668 24622
rect 45612 24518 45668 24556
rect 45612 23826 45668 23838
rect 45612 23774 45614 23826
rect 45666 23774 45668 23826
rect 44940 23266 45444 23268
rect 44940 23214 44942 23266
rect 44994 23214 45444 23266
rect 44940 23212 45444 23214
rect 44940 23202 44996 23212
rect 42812 23090 42868 23100
rect 42364 22146 42420 22158
rect 42364 22094 42366 22146
rect 42418 22094 42420 22146
rect 42028 21522 42084 21532
rect 42140 21700 42196 21710
rect 42364 21700 42420 22094
rect 42196 21644 42420 21700
rect 42140 21586 42196 21644
rect 42140 21534 42142 21586
rect 42194 21534 42196 21586
rect 42140 21522 42196 21534
rect 43484 21588 43540 21598
rect 42924 21476 42980 21486
rect 42924 21382 42980 21420
rect 41916 21308 42196 21364
rect 42140 20914 42196 21308
rect 42140 20862 42142 20914
rect 42194 20862 42196 20914
rect 42140 20850 42196 20862
rect 39900 19282 39956 19292
rect 40908 19348 40964 19358
rect 40908 19254 40964 19292
rect 41356 19348 41412 19358
rect 41468 19348 41524 20076
rect 42588 20578 42644 20590
rect 42588 20526 42590 20578
rect 42642 20526 42644 20578
rect 42588 20188 42644 20526
rect 43484 20356 43540 21532
rect 45052 21476 45108 21486
rect 45052 21382 45108 21420
rect 45388 20914 45444 23212
rect 45612 22372 45668 23774
rect 45612 21698 45668 22316
rect 45724 23826 45780 25788
rect 45724 23774 45726 23826
rect 45778 23774 45780 23826
rect 45724 22260 45780 23774
rect 45836 25618 45892 25630
rect 45836 25566 45838 25618
rect 45890 25566 45892 25618
rect 45836 24722 45892 25566
rect 45948 25506 46004 25788
rect 45948 25454 45950 25506
rect 46002 25454 46004 25506
rect 45948 25442 46004 25454
rect 46844 24948 46900 26126
rect 47516 26180 47572 26190
rect 47516 26086 47572 26124
rect 48076 25284 48132 26238
rect 48412 26292 48468 26302
rect 48524 26292 48580 26908
rect 48860 26404 48916 26414
rect 48412 26290 48580 26292
rect 48412 26238 48414 26290
rect 48466 26238 48580 26290
rect 48412 26236 48580 26238
rect 48748 26292 48804 26302
rect 48412 26226 48468 26236
rect 48748 26198 48804 26236
rect 48748 25508 48804 25518
rect 48748 25414 48804 25452
rect 48076 25218 48132 25228
rect 48412 25284 48468 25294
rect 48468 25228 48580 25284
rect 48412 25190 48468 25228
rect 46844 24882 46900 24892
rect 45836 24670 45838 24722
rect 45890 24670 45892 24722
rect 45836 23826 45892 24670
rect 47068 24052 47124 24062
rect 47068 23940 47124 23996
rect 45836 23774 45838 23826
rect 45890 23774 45892 23826
rect 45836 23380 45892 23774
rect 46956 23938 47124 23940
rect 46956 23886 47070 23938
rect 47122 23886 47124 23938
rect 46956 23884 47124 23886
rect 46284 23716 46340 23726
rect 46284 23714 46452 23716
rect 46284 23662 46286 23714
rect 46338 23662 46452 23714
rect 46284 23660 46452 23662
rect 46284 23650 46340 23660
rect 46396 23604 46452 23660
rect 46844 23714 46900 23726
rect 46844 23662 46846 23714
rect 46898 23662 46900 23714
rect 46844 23604 46900 23662
rect 46396 23538 46452 23548
rect 46508 23548 46900 23604
rect 46508 23380 46564 23548
rect 45836 23324 46564 23380
rect 46620 23380 46676 23390
rect 46172 22372 46228 22382
rect 45948 22370 46228 22372
rect 45948 22318 46174 22370
rect 46226 22318 46228 22370
rect 45948 22316 46228 22318
rect 45836 22260 45892 22270
rect 45724 22204 45836 22260
rect 45612 21646 45614 21698
rect 45666 21646 45668 21698
rect 45612 21476 45668 21646
rect 45836 21698 45892 22204
rect 45836 21646 45838 21698
rect 45890 21646 45892 21698
rect 45836 21634 45892 21646
rect 45612 21410 45668 21420
rect 45388 20862 45390 20914
rect 45442 20862 45444 20914
rect 45164 20804 45220 20814
rect 43484 20300 43988 20356
rect 42588 20132 42868 20188
rect 42588 20066 42644 20076
rect 41356 19346 41524 19348
rect 41356 19294 41358 19346
rect 41410 19294 41524 19346
rect 41356 19292 41524 19294
rect 41356 19236 41412 19292
rect 41356 19170 41412 19180
rect 38780 19122 38836 19134
rect 38780 19070 38782 19122
rect 38834 19070 38836 19122
rect 38780 18676 38836 19070
rect 38892 18676 38948 18686
rect 38780 18674 38948 18676
rect 38780 18622 38894 18674
rect 38946 18622 38948 18674
rect 38780 18620 38948 18622
rect 38892 18610 38948 18620
rect 37436 18398 37438 18450
rect 37490 18398 37492 18450
rect 37436 18386 37492 18398
rect 38220 18508 38612 18564
rect 36988 18286 36990 18338
rect 37042 18286 37044 18338
rect 36988 18274 37044 18286
rect 36764 17054 36766 17106
rect 36818 17054 36820 17106
rect 35196 16996 35252 17006
rect 34636 16830 34638 16882
rect 34690 16830 34692 16882
rect 34636 16818 34692 16830
rect 34860 16994 35252 16996
rect 34860 16942 35198 16994
rect 35250 16942 35252 16994
rect 34860 16940 35252 16942
rect 32956 16158 32958 16210
rect 33010 16158 33012 16210
rect 32956 16146 33012 16158
rect 30044 16100 30100 16110
rect 29932 16098 30100 16100
rect 29932 16046 30046 16098
rect 30098 16046 30100 16098
rect 29932 16044 30100 16046
rect 28028 13186 28196 13188
rect 28028 13134 28030 13186
rect 28082 13134 28196 13186
rect 28028 13132 28196 13134
rect 28252 13356 28644 13412
rect 29036 15202 29092 15214
rect 29036 15150 29038 15202
rect 29090 15150 29092 15202
rect 28252 13186 28308 13356
rect 28252 13134 28254 13186
rect 28306 13134 28308 13186
rect 28028 13122 28084 13132
rect 28252 13122 28308 13134
rect 28476 13188 28532 13198
rect 28476 13094 28532 13132
rect 29036 13188 29092 15150
rect 29036 13122 29092 13132
rect 29148 13634 29204 13646
rect 29148 13582 29150 13634
rect 29202 13582 29204 13634
rect 29148 13524 29204 13582
rect 28588 12850 28644 12862
rect 28588 12798 28590 12850
rect 28642 12798 28644 12850
rect 26348 12738 26404 12750
rect 26348 12686 26350 12738
rect 26402 12686 26404 12738
rect 26124 12066 26180 12078
rect 26124 12014 26126 12066
rect 26178 12014 26180 12066
rect 26124 11954 26180 12014
rect 26124 11902 26126 11954
rect 26178 11902 26180 11954
rect 26124 11620 26180 11902
rect 26124 11554 26180 11564
rect 26348 11508 26404 12686
rect 26684 12180 26740 12190
rect 26572 12178 26740 12180
rect 26572 12126 26686 12178
rect 26738 12126 26740 12178
rect 26572 12124 26740 12126
rect 26460 11956 26516 11966
rect 26572 11956 26628 12124
rect 26684 12114 26740 12124
rect 28028 12180 28084 12190
rect 28028 12086 28084 12124
rect 28588 12178 28644 12798
rect 28588 12126 28590 12178
rect 28642 12126 28644 12178
rect 28588 12114 28644 12126
rect 29148 12178 29204 13468
rect 29932 12964 29988 16044
rect 30044 16034 30100 16044
rect 33516 15876 33572 15886
rect 32732 15874 33572 15876
rect 32732 15822 33518 15874
rect 33570 15822 33572 15874
rect 32732 15820 33572 15822
rect 32732 14642 32788 15820
rect 33516 15810 33572 15820
rect 34076 15874 34132 15886
rect 34076 15822 34078 15874
rect 34130 15822 34132 15874
rect 32732 14590 32734 14642
rect 32786 14590 32788 14642
rect 32732 14578 32788 14590
rect 32060 14530 32116 14542
rect 32060 14478 32062 14530
rect 32114 14478 32116 14530
rect 29148 12126 29150 12178
rect 29202 12126 29204 12178
rect 29148 12114 29204 12126
rect 29820 12962 29988 12964
rect 29820 12910 29934 12962
rect 29986 12910 29988 12962
rect 29820 12908 29988 12910
rect 26460 11954 26628 11956
rect 26460 11902 26462 11954
rect 26514 11902 26628 11954
rect 26460 11900 26628 11902
rect 26684 11954 26740 11966
rect 26684 11902 26686 11954
rect 26738 11902 26740 11954
rect 26460 11890 26516 11900
rect 26348 11442 26404 11452
rect 25564 11342 25566 11394
rect 25618 11342 25620 11394
rect 25564 11330 25620 11342
rect 26236 11284 26292 11294
rect 26684 11284 26740 11902
rect 26236 11282 26740 11284
rect 26236 11230 26238 11282
rect 26290 11230 26740 11282
rect 26236 11228 26740 11230
rect 27020 11954 27076 11966
rect 27020 11902 27022 11954
rect 27074 11902 27076 11954
rect 26236 11218 26292 11228
rect 27020 10722 27076 11902
rect 28364 11956 28420 11966
rect 28364 11862 28420 11900
rect 29820 11844 29876 12908
rect 29932 12898 29988 12908
rect 30044 14306 30100 14318
rect 30940 14308 30996 14318
rect 30044 14254 30046 14306
rect 30098 14254 30100 14306
rect 29932 12292 29988 12302
rect 30044 12292 30100 14254
rect 30716 14306 30996 14308
rect 30716 14254 30942 14306
rect 30994 14254 30996 14306
rect 30716 14252 30996 14254
rect 30716 13074 30772 14252
rect 30940 14242 30996 14252
rect 32060 13972 32116 14478
rect 30716 13022 30718 13074
rect 30770 13022 30772 13074
rect 30716 13010 30772 13022
rect 31948 13916 32060 13972
rect 29932 12290 30100 12292
rect 29932 12238 29934 12290
rect 29986 12238 30100 12290
rect 29932 12236 30100 12238
rect 29932 12226 29988 12236
rect 28364 11506 28420 11518
rect 28364 11454 28366 11506
rect 28418 11454 28420 11506
rect 27020 10670 27022 10722
rect 27074 10670 27076 10722
rect 27020 10658 27076 10670
rect 27580 10668 27860 10724
rect 27580 10276 27636 10668
rect 27804 10612 27860 10668
rect 27916 10612 27972 10622
rect 28364 10612 28420 11454
rect 27804 10610 28420 10612
rect 27804 10558 27918 10610
rect 27970 10558 28420 10610
rect 27804 10556 28420 10558
rect 27916 10546 27972 10556
rect 27692 10500 27748 10510
rect 27692 10498 27860 10500
rect 27692 10446 27694 10498
rect 27746 10446 27860 10498
rect 27692 10444 27860 10446
rect 27692 10434 27748 10444
rect 27468 10220 27636 10276
rect 27804 10276 27860 10444
rect 27804 10220 27972 10276
rect 27468 9826 27524 10220
rect 27468 9774 27470 9826
rect 27522 9774 27524 9826
rect 27132 9714 27188 9726
rect 27132 9662 27134 9714
rect 27186 9662 27188 9714
rect 26908 9268 26964 9278
rect 26908 9174 26964 9212
rect 27132 9042 27188 9662
rect 27468 9154 27524 9774
rect 27580 9828 27636 9838
rect 27804 9828 27860 9838
rect 27916 9828 27972 10220
rect 27580 9734 27636 9772
rect 27692 9826 27972 9828
rect 27692 9774 27806 9826
rect 27858 9774 27972 9826
rect 27692 9772 27972 9774
rect 29820 9826 29876 11788
rect 31948 11844 32004 13916
rect 32060 13906 32116 13916
rect 33516 13972 33572 13982
rect 33516 13878 33572 13916
rect 34076 13972 34132 15822
rect 34860 14642 34916 16940
rect 35196 16930 35252 16940
rect 36764 16884 36820 17054
rect 37324 17108 37380 17118
rect 37324 16994 37380 17052
rect 37324 16942 37326 16994
rect 37378 16942 37380 16994
rect 37324 16930 37380 16942
rect 36764 16818 36820 16828
rect 37548 16884 37604 16894
rect 37548 16882 37716 16884
rect 37548 16830 37550 16882
rect 37602 16830 37716 16882
rect 37548 16828 37716 16830
rect 37548 16818 37604 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 37660 16322 37716 16828
rect 38220 16882 38276 18508
rect 40796 18452 40852 18462
rect 40796 18358 40852 18396
rect 41916 18452 41972 18462
rect 41916 18358 41972 18396
rect 41692 17666 41748 17678
rect 41692 17614 41694 17666
rect 41746 17614 41748 17666
rect 41020 17556 41076 17566
rect 41020 17462 41076 17500
rect 39788 16994 39844 17006
rect 39788 16942 39790 16994
rect 39842 16942 39844 16994
rect 38220 16830 38222 16882
rect 38274 16830 38276 16882
rect 38220 16818 38276 16830
rect 38556 16884 38612 16894
rect 38556 16790 38612 16828
rect 38556 16658 38612 16670
rect 38556 16606 38558 16658
rect 38610 16606 38612 16658
rect 37660 16270 37662 16322
rect 37714 16270 37716 16322
rect 37660 16258 37716 16270
rect 37996 16324 38052 16334
rect 37996 16322 38500 16324
rect 37996 16270 37998 16322
rect 38050 16270 38500 16322
rect 37996 16268 38500 16270
rect 37996 16258 38052 16268
rect 37772 16212 37828 16222
rect 37772 16118 37828 16156
rect 38220 16098 38276 16110
rect 38220 16046 38222 16098
rect 38274 16046 38276 16098
rect 36428 15874 36484 15886
rect 36428 15822 36430 15874
rect 36482 15822 36484 15874
rect 36316 15428 36372 15438
rect 36428 15428 36484 15822
rect 36316 15426 36484 15428
rect 36316 15374 36318 15426
rect 36370 15374 36484 15426
rect 36316 15372 36484 15374
rect 36316 15362 36372 15372
rect 35644 15314 35700 15326
rect 35644 15262 35646 15314
rect 35698 15262 35700 15314
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34860 14590 34862 14642
rect 34914 14590 34916 14642
rect 34860 14578 34916 14590
rect 34076 13906 34132 13916
rect 35308 14306 35364 14318
rect 35308 14254 35310 14306
rect 35362 14254 35364 14306
rect 35308 13972 35364 14254
rect 35308 13906 35364 13916
rect 35532 13748 35588 13758
rect 35644 13748 35700 15262
rect 36316 14306 36372 14318
rect 36316 14254 36318 14306
rect 36370 14254 36372 14306
rect 36204 13860 36260 13870
rect 36316 13860 36372 14254
rect 36204 13858 36372 13860
rect 36204 13806 36206 13858
rect 36258 13806 36372 13858
rect 36204 13804 36372 13806
rect 36204 13794 36260 13804
rect 35532 13746 35700 13748
rect 35532 13694 35534 13746
rect 35586 13694 35700 13746
rect 35532 13692 35700 13694
rect 35532 13682 35588 13692
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 32844 13076 32900 13086
rect 33404 13076 33460 13086
rect 32508 13074 32900 13076
rect 32508 13022 32846 13074
rect 32898 13022 32900 13074
rect 32508 13020 32900 13022
rect 31948 11506 32004 11788
rect 31948 11454 31950 11506
rect 32002 11454 32004 11506
rect 31948 9940 32004 11454
rect 32060 12066 32116 12078
rect 32060 12014 32062 12066
rect 32114 12014 32116 12066
rect 32060 10612 32116 12014
rect 32172 11956 32228 11966
rect 32172 10834 32228 11900
rect 32172 10782 32174 10834
rect 32226 10782 32228 10834
rect 32172 10770 32228 10782
rect 32284 10612 32340 10622
rect 32060 10610 32340 10612
rect 32060 10558 32286 10610
rect 32338 10558 32340 10610
rect 32060 10556 32340 10558
rect 32284 10546 32340 10556
rect 32508 10610 32564 13020
rect 32844 13010 32900 13020
rect 32956 13074 33460 13076
rect 32956 13022 33406 13074
rect 33458 13022 33460 13074
rect 32956 13020 33460 13022
rect 32508 10558 32510 10610
rect 32562 10558 32564 10610
rect 32508 10546 32564 10558
rect 32732 10612 32788 10622
rect 32956 10612 33012 13020
rect 33404 13010 33460 13020
rect 35644 12964 35700 13692
rect 38220 13636 38276 16046
rect 38444 15202 38500 16268
rect 38444 15150 38446 15202
rect 38498 15150 38500 15202
rect 38444 15138 38500 15150
rect 38332 13636 38388 13646
rect 38220 13634 38388 13636
rect 38220 13582 38334 13634
rect 38386 13582 38388 13634
rect 38220 13580 38388 13582
rect 38332 13570 38388 13580
rect 35644 12898 35700 12908
rect 36316 12964 36372 12974
rect 35532 12850 35588 12862
rect 35532 12798 35534 12850
rect 35586 12798 35588 12850
rect 33964 12404 34020 12414
rect 33964 12310 34020 12348
rect 35532 12404 35588 12798
rect 36316 12740 36372 12908
rect 36764 12740 36820 12750
rect 36316 12738 36820 12740
rect 36316 12686 36766 12738
rect 36818 12686 36820 12738
rect 36316 12684 36820 12686
rect 36764 12404 36820 12684
rect 36988 12404 37044 12414
rect 36764 12348 36988 12404
rect 35532 12338 35588 12348
rect 36988 12178 37044 12348
rect 36988 12126 36990 12178
rect 37042 12126 37044 12178
rect 36988 12114 37044 12126
rect 37660 12068 37716 12078
rect 37660 12066 38500 12068
rect 37660 12014 37662 12066
rect 37714 12014 38500 12066
rect 37660 12012 38500 12014
rect 37660 12002 37716 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 38332 11620 38388 11630
rect 35756 11508 35812 11518
rect 35756 11394 35812 11452
rect 36204 11508 36260 11518
rect 36204 11414 36260 11452
rect 35756 11342 35758 11394
rect 35810 11342 35812 11394
rect 35756 11330 35812 11342
rect 32732 10610 33012 10612
rect 32732 10558 32734 10610
rect 32786 10558 33012 10610
rect 32732 10556 33012 10558
rect 38332 10612 38388 11564
rect 38444 11506 38500 12012
rect 38556 11620 38612 16606
rect 38780 16212 38836 16222
rect 38780 16118 38836 16156
rect 39788 16212 39844 16942
rect 39788 16146 39844 16156
rect 40908 16212 40964 16222
rect 40908 16118 40964 16156
rect 41692 16098 41748 17614
rect 42364 17556 42420 17566
rect 42364 17462 42420 17500
rect 42812 16884 42868 20132
rect 43708 20130 43764 20142
rect 43708 20078 43710 20130
rect 43762 20078 43764 20130
rect 43708 18452 43764 20078
rect 43932 20132 43988 20300
rect 43932 18562 43988 20076
rect 45164 19906 45220 20748
rect 45388 20188 45444 20862
rect 45948 20804 46004 22316
rect 46172 22306 46228 22316
rect 46284 22372 46340 22382
rect 46284 22258 46340 22316
rect 46284 22206 46286 22258
rect 46338 22206 46340 22258
rect 46284 22194 46340 22206
rect 46060 21924 46116 21934
rect 46396 21924 46452 23324
rect 46508 22260 46564 22270
rect 46508 22166 46564 22204
rect 46060 21810 46116 21868
rect 46060 21758 46062 21810
rect 46114 21758 46116 21810
rect 46060 21746 46116 21758
rect 46284 21868 46452 21924
rect 46284 21586 46340 21868
rect 46284 21534 46286 21586
rect 46338 21534 46340 21586
rect 46284 21522 46340 21534
rect 46396 21698 46452 21710
rect 46396 21646 46398 21698
rect 46450 21646 46452 21698
rect 46172 20916 46228 20926
rect 46396 20916 46452 21646
rect 46172 20914 46452 20916
rect 46172 20862 46174 20914
rect 46226 20862 46452 20914
rect 46172 20860 46452 20862
rect 46172 20850 46228 20860
rect 45948 20672 46004 20748
rect 46284 20692 46340 20702
rect 46620 20692 46676 23324
rect 46956 22370 47012 23884
rect 47068 23874 47124 23884
rect 48300 23938 48356 23950
rect 48300 23886 48302 23938
rect 48354 23886 48356 23938
rect 47964 23716 48020 23726
rect 47740 23492 47796 23502
rect 47292 23042 47348 23054
rect 47292 22990 47294 23042
rect 47346 22990 47348 23042
rect 47180 22596 47236 22606
rect 47180 22502 47236 22540
rect 46956 22318 46958 22370
rect 47010 22318 47012 22370
rect 46956 22306 47012 22318
rect 47068 22372 47124 22382
rect 47292 22372 47348 22990
rect 46844 21698 46900 21710
rect 46844 21646 46846 21698
rect 46898 21646 46900 21698
rect 46844 21586 46900 21646
rect 46844 21534 46846 21586
rect 46898 21534 46900 21586
rect 46844 21522 46900 21534
rect 47068 21586 47124 22316
rect 47068 21534 47070 21586
rect 47122 21534 47124 21586
rect 47068 21522 47124 21534
rect 47180 22316 47348 22372
rect 47404 22708 47460 22718
rect 47180 21924 47236 22316
rect 46284 20690 46676 20692
rect 46284 20638 46286 20690
rect 46338 20638 46676 20690
rect 46284 20636 46676 20638
rect 46284 20626 46340 20636
rect 45388 20132 45556 20188
rect 45164 19854 45166 19906
rect 45218 19854 45220 19906
rect 45164 19842 45220 19854
rect 43932 18510 43934 18562
rect 43986 18510 43988 18562
rect 43932 18498 43988 18510
rect 43484 18396 43764 18452
rect 43484 16994 43540 18396
rect 45500 18116 45556 20132
rect 47180 20132 47236 21868
rect 47292 21588 47348 21598
rect 47404 21588 47460 22652
rect 47740 22594 47796 23436
rect 47740 22542 47742 22594
rect 47794 22542 47796 22594
rect 47740 22530 47796 22542
rect 47964 22372 48020 23660
rect 48076 23714 48132 23726
rect 48076 23662 48078 23714
rect 48130 23662 48132 23714
rect 48076 23380 48132 23662
rect 48076 22708 48132 23324
rect 48076 22642 48132 22652
rect 48300 23156 48356 23886
rect 48524 23378 48580 25228
rect 48860 24946 48916 26348
rect 49420 25172 49476 27804
rect 49532 27794 49588 27804
rect 49756 27860 49812 28590
rect 49756 27794 49812 27804
rect 49868 27074 49924 27086
rect 50092 27076 50148 29150
rect 52668 28754 52724 28766
rect 52668 28702 52670 28754
rect 52722 28702 52724 28754
rect 50540 28532 50596 28542
rect 50540 28530 51380 28532
rect 50540 28478 50542 28530
rect 50594 28478 51380 28530
rect 50540 28476 51380 28478
rect 50540 28466 50596 28476
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 49868 27022 49870 27074
rect 49922 27022 49924 27074
rect 49756 26964 49812 26974
rect 49868 26964 49924 27022
rect 49812 26908 49924 26964
rect 49980 27074 50148 27076
rect 49980 27022 50094 27074
rect 50146 27022 50148 27074
rect 49980 27020 50148 27022
rect 49756 26514 49812 26908
rect 49756 26462 49758 26514
rect 49810 26462 49812 26514
rect 49756 26450 49812 26462
rect 49644 26404 49700 26414
rect 49532 26292 49588 26302
rect 49532 25396 49588 26236
rect 49644 25620 49700 26348
rect 49868 26404 49924 26442
rect 49868 26338 49924 26348
rect 49980 26402 50036 27020
rect 50092 27010 50148 27020
rect 50204 27076 50260 27086
rect 50204 27074 50484 27076
rect 50204 27022 50206 27074
rect 50258 27022 50484 27074
rect 50204 27020 50484 27022
rect 50204 27010 50260 27020
rect 49980 26350 49982 26402
rect 50034 26350 50036 26402
rect 49644 25508 49700 25564
rect 49868 26178 49924 26190
rect 49868 26126 49870 26178
rect 49922 26126 49924 26178
rect 49756 25508 49812 25518
rect 49644 25506 49812 25508
rect 49644 25454 49758 25506
rect 49810 25454 49812 25506
rect 49644 25452 49812 25454
rect 49756 25442 49812 25452
rect 49868 25508 49924 26126
rect 49532 25302 49588 25340
rect 49420 25116 49700 25172
rect 48860 24894 48862 24946
rect 48914 24894 48916 24946
rect 48860 24882 48916 24894
rect 49532 24834 49588 24846
rect 49532 24782 49534 24834
rect 49586 24782 49588 24834
rect 49532 23716 49588 24782
rect 49532 23650 49588 23660
rect 48524 23326 48526 23378
rect 48578 23326 48580 23378
rect 48524 23314 48580 23326
rect 48300 22596 48356 23100
rect 48748 23156 48804 23166
rect 49532 23156 49588 23166
rect 48748 23154 49588 23156
rect 48748 23102 48750 23154
rect 48802 23102 49534 23154
rect 49586 23102 49588 23154
rect 48748 23100 49588 23102
rect 48748 23090 48804 23100
rect 49532 23090 49588 23100
rect 48300 22530 48356 22540
rect 48636 23042 48692 23054
rect 48636 22990 48638 23042
rect 48690 22990 48692 23042
rect 47964 22278 48020 22316
rect 48076 22370 48132 22382
rect 48076 22318 48078 22370
rect 48130 22318 48132 22370
rect 47292 21586 47460 21588
rect 47292 21534 47294 21586
rect 47346 21534 47460 21586
rect 47292 21532 47460 21534
rect 47628 22258 47684 22270
rect 47628 22206 47630 22258
rect 47682 22206 47684 22258
rect 47628 21588 47684 22206
rect 48076 22036 48132 22318
rect 48076 21970 48132 21980
rect 47292 21522 47348 21532
rect 47628 21522 47684 21532
rect 47404 21362 47460 21374
rect 47404 21310 47406 21362
rect 47458 21310 47460 21362
rect 45388 18060 45556 18116
rect 46508 19010 46564 19022
rect 46508 18958 46510 19010
rect 46562 18958 46564 19010
rect 43484 16942 43486 16994
rect 43538 16942 43540 16994
rect 43484 16930 43540 16942
rect 44492 17778 44548 17790
rect 44492 17726 44494 17778
rect 44546 17726 44548 17778
rect 42812 16790 42868 16828
rect 41692 16046 41694 16098
rect 41746 16046 41748 16098
rect 38892 15876 38948 15886
rect 38892 15538 38948 15820
rect 38892 15486 38894 15538
rect 38946 15486 38948 15538
rect 38780 13972 38836 13982
rect 38892 13972 38948 15486
rect 41692 15876 41748 16046
rect 44044 15988 44100 15998
rect 44044 15894 44100 15932
rect 38780 13970 38948 13972
rect 38780 13918 38782 13970
rect 38834 13918 38948 13970
rect 38780 13916 38948 13918
rect 38780 13906 38836 13916
rect 38892 12404 38948 13916
rect 39564 14644 39620 14654
rect 39564 14530 39620 14588
rect 41692 14642 41748 15820
rect 42140 15876 42196 15886
rect 42140 15782 42196 15820
rect 41692 14590 41694 14642
rect 41746 14590 41748 14642
rect 41692 14578 41748 14590
rect 42252 15426 42308 15438
rect 42252 15374 42254 15426
rect 42306 15374 42308 15426
rect 39564 14478 39566 14530
rect 39618 14478 39620 14530
rect 39116 12964 39172 12974
rect 39116 12870 39172 12908
rect 38892 12338 38948 12348
rect 38556 11554 38612 11564
rect 39116 11620 39172 11630
rect 38444 11454 38446 11506
rect 38498 11454 38500 11506
rect 38444 11442 38500 11454
rect 39116 11506 39172 11564
rect 39116 11454 39118 11506
rect 39170 11454 39172 11506
rect 39116 11442 39172 11454
rect 39564 11508 39620 14478
rect 40012 13860 40068 13870
rect 39788 13858 40068 13860
rect 39788 13806 40014 13858
rect 40066 13806 40068 13858
rect 39788 13804 40068 13806
rect 39788 13074 39844 13804
rect 40012 13794 40068 13804
rect 39788 13022 39790 13074
rect 39842 13022 39844 13074
rect 39788 13010 39844 13022
rect 41916 13076 41972 13086
rect 41916 12982 41972 13020
rect 41580 12964 41636 12974
rect 40236 12404 40292 12414
rect 40236 12310 40292 12348
rect 41580 12180 41636 12908
rect 42252 12292 42308 15374
rect 44492 15316 44548 17726
rect 45388 16884 45444 18060
rect 45500 17780 45556 17790
rect 46508 17780 46564 18958
rect 45500 17778 46340 17780
rect 45500 17726 45502 17778
rect 45554 17726 46340 17778
rect 45500 17724 46340 17726
rect 45500 17714 45556 17724
rect 45388 16818 45444 16828
rect 46060 16884 46116 16894
rect 46060 16790 46116 16828
rect 45612 16772 45668 16782
rect 45612 16770 46004 16772
rect 45612 16718 45614 16770
rect 45666 16718 46004 16770
rect 45612 16716 46004 16718
rect 45612 16706 45668 16716
rect 45500 16212 45556 16222
rect 45500 16210 45892 16212
rect 45500 16158 45502 16210
rect 45554 16158 45892 16210
rect 45500 16156 45892 16158
rect 45500 16146 45556 16156
rect 44716 15876 44772 15886
rect 44716 15782 44772 15820
rect 44492 15250 44548 15260
rect 45612 15316 45668 15326
rect 45612 15222 45668 15260
rect 45836 15314 45892 16156
rect 45836 15262 45838 15314
rect 45890 15262 45892 15314
rect 45836 15250 45892 15262
rect 45948 15316 46004 16716
rect 46060 15316 46116 15326
rect 45948 15314 46116 15316
rect 45948 15262 46062 15314
rect 46114 15262 46116 15314
rect 45948 15260 46116 15262
rect 46060 15250 46116 15260
rect 46284 15314 46340 17724
rect 46508 17714 46564 17724
rect 47180 17108 47236 20076
rect 47292 20132 47348 20142
rect 47404 20132 47460 21310
rect 48636 20916 48692 22990
rect 49644 21924 49700 25116
rect 49868 24834 49924 25452
rect 49980 25394 50036 26350
rect 50204 26740 50260 26750
rect 50092 25732 50148 25742
rect 50204 25732 50260 26684
rect 50092 25730 50260 25732
rect 50092 25678 50094 25730
rect 50146 25678 50260 25730
rect 50092 25676 50260 25678
rect 50092 25666 50148 25676
rect 50428 25620 50484 27020
rect 51212 26962 51268 26974
rect 51212 26910 51214 26962
rect 51266 26910 51268 26962
rect 50652 26852 50708 26890
rect 50652 26786 50708 26796
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50428 25526 50484 25564
rect 50988 26404 51044 26414
rect 49980 25342 49982 25394
rect 50034 25342 50036 25394
rect 49980 25330 50036 25342
rect 50876 25396 50932 25406
rect 50876 25302 50932 25340
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 49868 24782 49870 24834
rect 49922 24782 49924 24834
rect 49868 24770 49924 24782
rect 50988 24948 51044 26348
rect 51100 26292 51156 26302
rect 51100 25506 51156 26236
rect 51212 25620 51268 26910
rect 51324 26850 51380 28476
rect 52108 27860 52164 27870
rect 52108 27746 52164 27804
rect 52108 27694 52110 27746
rect 52162 27694 52164 27746
rect 52108 27682 52164 27694
rect 52444 27188 52500 27198
rect 52668 27188 52724 28702
rect 52444 27186 52724 27188
rect 52444 27134 52446 27186
rect 52498 27134 52724 27186
rect 52444 27132 52724 27134
rect 53340 28418 53396 28430
rect 53340 28366 53342 28418
rect 53394 28366 53396 28418
rect 53340 27860 53396 28366
rect 51660 27076 51716 27086
rect 51548 26964 51604 27002
rect 51660 26982 51716 27020
rect 51548 26898 51604 26908
rect 52332 26964 52388 27002
rect 52332 26898 52388 26908
rect 51324 26798 51326 26850
rect 51378 26798 51380 26850
rect 51324 26786 51380 26798
rect 51324 26404 51380 26414
rect 51324 26310 51380 26348
rect 51436 26292 51492 26302
rect 51492 26236 51716 26292
rect 51436 26198 51492 26236
rect 51324 26068 51380 26078
rect 51324 26066 51492 26068
rect 51324 26014 51326 26066
rect 51378 26014 51492 26066
rect 51324 26012 51492 26014
rect 51324 26002 51380 26012
rect 51212 25564 51380 25620
rect 51100 25454 51102 25506
rect 51154 25454 51156 25506
rect 51100 25442 51156 25454
rect 51212 25394 51268 25406
rect 51212 25342 51214 25394
rect 51266 25342 51268 25394
rect 51212 24948 51268 25342
rect 50988 24892 51268 24948
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 49756 23156 49812 23166
rect 49756 23062 49812 23100
rect 50428 23154 50484 23166
rect 50428 23102 50430 23154
rect 50482 23102 50484 23154
rect 49644 21858 49700 21868
rect 50428 22932 50484 23102
rect 50988 23156 51044 24892
rect 51212 24724 51268 24734
rect 51100 24668 51212 24724
rect 51100 23826 51156 24668
rect 51212 24592 51268 24668
rect 51324 24050 51380 25564
rect 51436 24610 51492 26012
rect 51548 25506 51604 25518
rect 51548 25454 51550 25506
rect 51602 25454 51604 25506
rect 51548 24724 51604 25454
rect 51548 24658 51604 24668
rect 51436 24558 51438 24610
rect 51490 24558 51492 24610
rect 51436 24546 51492 24558
rect 51324 23998 51326 24050
rect 51378 23998 51380 24050
rect 51324 23986 51380 23998
rect 51660 23940 51716 26236
rect 52444 25506 52500 27132
rect 53340 27076 53396 27804
rect 56700 27186 56756 27198
rect 56700 27134 56702 27186
rect 56754 27134 56756 27186
rect 53788 27076 53844 27086
rect 53340 27074 53844 27076
rect 53340 27022 53790 27074
rect 53842 27022 53844 27074
rect 53340 27020 53844 27022
rect 53228 26516 53284 26526
rect 53340 26516 53396 27020
rect 53788 27010 53844 27020
rect 54572 26962 54628 26974
rect 54572 26910 54574 26962
rect 54626 26910 54628 26962
rect 54572 26908 54628 26910
rect 53228 26514 53396 26516
rect 53228 26462 53230 26514
rect 53282 26462 53396 26514
rect 53228 26460 53396 26462
rect 53676 26852 53732 26862
rect 53228 26450 53284 26460
rect 53676 26402 53732 26796
rect 54012 26852 54628 26908
rect 55356 26964 55412 26974
rect 54012 26514 54068 26852
rect 54012 26462 54014 26514
rect 54066 26462 54068 26514
rect 54012 26450 54068 26462
rect 53676 26350 53678 26402
rect 53730 26350 53732 26402
rect 53676 26338 53732 26350
rect 55356 26178 55412 26908
rect 56140 26292 56196 26302
rect 56700 26292 56756 27134
rect 56140 26290 56756 26292
rect 56140 26238 56142 26290
rect 56194 26238 56756 26290
rect 56140 26236 56756 26238
rect 56140 26226 56196 26236
rect 55356 26126 55358 26178
rect 55410 26126 55412 26178
rect 55356 26114 55412 26126
rect 52444 25454 52446 25506
rect 52498 25454 52500 25506
rect 52444 25442 52500 25454
rect 52444 24724 52500 24734
rect 51884 24612 51940 24622
rect 51884 24610 52388 24612
rect 51884 24558 51886 24610
rect 51938 24558 52388 24610
rect 51884 24556 52388 24558
rect 51884 24546 51940 24556
rect 52332 24162 52388 24556
rect 52444 24610 52500 24668
rect 55356 24722 55412 24734
rect 55356 24670 55358 24722
rect 55410 24670 55412 24722
rect 52444 24558 52446 24610
rect 52498 24558 52500 24610
rect 52444 24546 52500 24558
rect 54572 24610 54628 24622
rect 54572 24558 54574 24610
rect 54626 24558 54628 24610
rect 52332 24110 52334 24162
rect 52386 24110 52388 24162
rect 52332 24098 52388 24110
rect 52668 24164 52724 24174
rect 52668 24070 52724 24108
rect 54572 24164 54628 24558
rect 54572 24098 54628 24108
rect 55356 24612 55412 24670
rect 51100 23774 51102 23826
rect 51154 23774 51156 23826
rect 51100 23762 51156 23774
rect 51436 23938 51716 23940
rect 51436 23886 51662 23938
rect 51714 23886 51716 23938
rect 51436 23884 51716 23886
rect 51324 23714 51380 23726
rect 51324 23662 51326 23714
rect 51378 23662 51380 23714
rect 51324 23604 51380 23662
rect 50988 23090 51044 23100
rect 51100 23548 51380 23604
rect 51100 23380 51156 23548
rect 48748 20916 48804 20926
rect 48636 20914 48804 20916
rect 48636 20862 48750 20914
rect 48802 20862 48804 20914
rect 48636 20860 48804 20862
rect 50428 20916 50484 22876
rect 51100 22372 51156 23324
rect 51100 22306 51156 22316
rect 51212 23380 51268 23390
rect 51436 23380 51492 23884
rect 51660 23874 51716 23884
rect 51212 23378 51492 23380
rect 51212 23326 51214 23378
rect 51266 23326 51492 23378
rect 51212 23324 51492 23326
rect 51660 23716 51716 23726
rect 51212 22370 51268 23324
rect 51548 22932 51604 22942
rect 51548 22838 51604 22876
rect 51660 22594 51716 23660
rect 52556 23716 52612 23726
rect 52556 23622 52612 23660
rect 52220 23380 52276 23390
rect 51660 22542 51662 22594
rect 51714 22542 51716 22594
rect 51660 22530 51716 22542
rect 51772 23156 51828 23166
rect 51772 23042 51828 23100
rect 52220 23154 52276 23324
rect 52220 23102 52222 23154
rect 52274 23102 52276 23154
rect 52220 23090 52276 23102
rect 52556 23154 52612 23166
rect 52556 23102 52558 23154
rect 52610 23102 52612 23154
rect 51772 22990 51774 23042
rect 51826 22990 51828 23042
rect 51212 22318 51214 22370
rect 51266 22318 51268 22370
rect 51212 22306 51268 22318
rect 51436 22372 51492 22382
rect 51436 22278 51492 22316
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50876 21812 50932 21822
rect 50876 21718 50932 21756
rect 51436 21812 51492 21822
rect 51436 21586 51492 21756
rect 51436 21534 51438 21586
rect 51490 21534 51492 21586
rect 51436 21522 51492 21534
rect 50876 20916 50932 20926
rect 50428 20914 50932 20916
rect 50428 20862 50878 20914
rect 50930 20862 50932 20914
rect 50428 20860 50932 20862
rect 48748 20850 48804 20860
rect 50876 20850 50932 20860
rect 47292 20130 47460 20132
rect 47292 20078 47294 20130
rect 47346 20078 47460 20130
rect 47292 20076 47460 20078
rect 48076 20802 48132 20814
rect 48076 20750 48078 20802
rect 48130 20750 48132 20802
rect 47292 20066 47348 20076
rect 48076 20018 48132 20750
rect 51324 20578 51380 20590
rect 51324 20526 51326 20578
rect 51378 20526 51380 20578
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 48076 19966 48078 20018
rect 48130 19966 48132 20018
rect 48076 19908 48132 19966
rect 49644 20244 49700 20254
rect 48524 19908 48580 19918
rect 48076 19906 48580 19908
rect 48076 19854 48526 19906
rect 48578 19854 48580 19906
rect 48076 19852 48580 19854
rect 48524 19236 48580 19852
rect 49644 19346 49700 20188
rect 50540 20244 50596 20282
rect 50540 20178 50596 20188
rect 49980 20132 50036 20142
rect 49980 20130 50372 20132
rect 49980 20078 49982 20130
rect 50034 20078 50372 20130
rect 49980 20076 50372 20078
rect 49980 20066 50036 20076
rect 49644 19294 49646 19346
rect 49698 19294 49700 19346
rect 49644 19282 49700 19294
rect 48860 19236 48916 19246
rect 48524 19234 48916 19236
rect 48524 19182 48862 19234
rect 48914 19182 48916 19234
rect 48524 19180 48916 19182
rect 47628 17780 47684 17790
rect 47628 17686 47684 17724
rect 46284 15262 46286 15314
rect 46338 15262 46340 15314
rect 46284 15250 46340 15262
rect 46956 17052 47180 17108
rect 46396 15092 46452 15102
rect 46396 15090 46900 15092
rect 46396 15038 46398 15090
rect 46450 15038 46900 15090
rect 46396 15036 46900 15038
rect 46396 15026 46452 15036
rect 43820 14644 43876 14654
rect 43820 14550 43876 14588
rect 46284 14306 46340 14318
rect 46284 14254 46286 14306
rect 46338 14254 46340 14306
rect 45388 13634 45444 13646
rect 45388 13582 45390 13634
rect 45442 13582 45444 13634
rect 45388 12964 45444 13582
rect 45836 13076 45892 13086
rect 45500 12964 45556 12974
rect 45388 12962 45556 12964
rect 45388 12910 45502 12962
rect 45554 12910 45556 12962
rect 45388 12908 45556 12910
rect 44044 12852 44100 12862
rect 44044 12758 44100 12796
rect 42364 12292 42420 12302
rect 42252 12290 42420 12292
rect 42252 12238 42366 12290
rect 42418 12238 42420 12290
rect 42252 12236 42420 12238
rect 42364 12226 42420 12236
rect 39564 11442 39620 11452
rect 39788 12066 39844 12078
rect 39788 12014 39790 12066
rect 39842 12014 39844 12066
rect 41580 12048 41636 12124
rect 45276 12180 45332 12190
rect 45388 12180 45444 12908
rect 45500 12898 45556 12908
rect 45332 12124 45444 12180
rect 45276 12114 45332 12124
rect 44492 12066 44548 12078
rect 38556 11172 38612 11182
rect 38556 11078 38612 11116
rect 39228 11172 39284 11182
rect 38444 10612 38500 10622
rect 38332 10610 38500 10612
rect 38332 10558 38446 10610
rect 38498 10558 38500 10610
rect 38332 10556 38500 10558
rect 32732 10546 32788 10556
rect 32172 10386 32228 10398
rect 32172 10334 32174 10386
rect 32226 10334 32228 10386
rect 32172 10164 32228 10334
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 32172 10108 32676 10164
rect 35196 10154 35460 10164
rect 38332 10164 38388 10556
rect 38444 10546 38500 10556
rect 39228 10612 39284 11116
rect 39788 11172 39844 12014
rect 44492 12014 44494 12066
rect 44546 12014 44548 12066
rect 39788 11106 39844 11116
rect 40012 11620 40068 11630
rect 40012 10834 40068 11564
rect 44492 11620 44548 12014
rect 45500 12068 45556 12078
rect 45500 12066 45668 12068
rect 45500 12014 45502 12066
rect 45554 12014 45668 12066
rect 45500 12012 45668 12014
rect 45500 12002 45556 12012
rect 44492 11554 44548 11564
rect 45612 11396 45668 12012
rect 45724 11620 45780 11630
rect 45724 11526 45780 11564
rect 45836 11618 45892 13020
rect 46284 13076 46340 14254
rect 46284 13010 46340 13020
rect 46284 12852 46340 12862
rect 46284 12758 46340 12796
rect 46396 12404 46452 12414
rect 45836 11566 45838 11618
rect 45890 11566 45892 11618
rect 45836 11554 45892 11566
rect 46060 11844 46116 11854
rect 46060 11618 46116 11788
rect 46396 11844 46452 12348
rect 46396 11778 46452 11788
rect 46060 11566 46062 11618
rect 46114 11566 46116 11618
rect 46060 11554 46116 11566
rect 46284 11396 46340 11406
rect 45612 11394 46340 11396
rect 45612 11342 46286 11394
rect 46338 11342 46340 11394
rect 45612 11340 46340 11342
rect 46284 11330 46340 11340
rect 46844 11394 46900 15036
rect 46956 14644 47012 17052
rect 47180 17042 47236 17052
rect 48300 17666 48356 17678
rect 48300 17614 48302 17666
rect 48354 17614 48356 17666
rect 48300 17444 48356 17614
rect 48300 16770 48356 17388
rect 48860 17444 48916 19180
rect 48860 17350 48916 17388
rect 49644 18452 49700 18462
rect 49644 17444 49700 18396
rect 50316 18450 50372 20076
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50316 18398 50318 18450
rect 50370 18398 50372 18450
rect 50316 18386 50372 18398
rect 51324 18452 51380 20526
rect 51772 20188 51828 22990
rect 52444 23042 52500 23054
rect 52444 22990 52446 23042
rect 52498 22990 52500 23042
rect 52444 22708 52500 22990
rect 52556 22932 52612 23102
rect 52780 23156 52836 23166
rect 52780 23062 52836 23100
rect 52556 22866 52612 22876
rect 51996 22652 52500 22708
rect 51996 22370 52052 22652
rect 51996 22318 51998 22370
rect 52050 22318 52052 22370
rect 51996 22306 52052 22318
rect 51996 22146 52052 22158
rect 51996 22094 51998 22146
rect 52050 22094 52052 22146
rect 51996 21252 52052 22094
rect 55356 21700 55412 24556
rect 55916 24612 55972 24622
rect 55916 24518 55972 24556
rect 54908 21698 55412 21700
rect 54908 21646 55358 21698
rect 55410 21646 55412 21698
rect 54908 21644 55412 21646
rect 51996 21186 52052 21196
rect 53676 21252 53732 21262
rect 51548 20132 51828 20188
rect 51548 19906 51604 20132
rect 53676 20130 53732 21196
rect 53676 20078 53678 20130
rect 53730 20078 53732 20130
rect 53676 20066 53732 20078
rect 54908 20242 54964 21644
rect 55356 21634 55412 21644
rect 54908 20190 54910 20242
rect 54962 20190 54964 20242
rect 54460 20020 54516 20030
rect 54908 20020 54964 20190
rect 54460 20018 54964 20020
rect 54460 19966 54462 20018
rect 54514 19966 54964 20018
rect 54460 19964 54964 19966
rect 54460 19954 54516 19964
rect 51548 19854 51550 19906
rect 51602 19854 51604 19906
rect 51548 19842 51604 19854
rect 51772 19346 51828 19358
rect 51772 19294 51774 19346
rect 51826 19294 51828 19346
rect 51380 18396 51604 18452
rect 51324 18386 51380 18396
rect 48748 17108 48804 17118
rect 48748 17014 48804 17052
rect 49532 17108 49588 17118
rect 49532 16882 49588 17052
rect 49532 16830 49534 16882
rect 49586 16830 49588 16882
rect 49532 16818 49588 16830
rect 48300 16718 48302 16770
rect 48354 16718 48356 16770
rect 48300 16098 48356 16718
rect 48300 16046 48302 16098
rect 48354 16046 48356 16098
rect 47628 15988 47684 15998
rect 47628 15894 47684 15932
rect 48300 15764 48356 16046
rect 49644 16100 49700 17388
rect 51548 17444 51604 18396
rect 51772 18228 51828 19294
rect 53452 19346 53508 19358
rect 53452 19294 53454 19346
rect 53506 19294 53508 19346
rect 52668 19124 52724 19134
rect 52668 19030 52724 19068
rect 53340 18452 53396 18462
rect 52444 18450 53396 18452
rect 52444 18398 53342 18450
rect 53394 18398 53396 18450
rect 52444 18396 53396 18398
rect 53452 18452 53508 19294
rect 54908 19236 54964 19964
rect 54908 19170 54964 19180
rect 56252 19236 56308 19246
rect 56252 19142 56308 19180
rect 56812 19236 56868 19246
rect 55580 19124 55636 19134
rect 55580 19030 55636 19068
rect 53676 18674 53732 18686
rect 53676 18622 53678 18674
rect 53730 18622 53732 18674
rect 53564 18452 53620 18462
rect 53452 18450 53620 18452
rect 53452 18398 53566 18450
rect 53618 18398 53620 18450
rect 53452 18396 53620 18398
rect 52444 18338 52500 18396
rect 53340 18386 53396 18396
rect 53564 18386 53620 18396
rect 52444 18286 52446 18338
rect 52498 18286 52500 18338
rect 52444 18274 52500 18286
rect 51772 18162 51828 18172
rect 53228 18228 53284 18238
rect 53228 18134 53284 18172
rect 51996 17444 52052 17454
rect 51548 17388 51996 17444
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 51548 16994 51604 17388
rect 51996 17312 52052 17388
rect 52668 17444 52724 17454
rect 52724 17388 52948 17444
rect 52668 17350 52724 17388
rect 51548 16942 51550 16994
rect 51602 16942 51604 16994
rect 51548 16930 51604 16942
rect 52668 16212 52724 16222
rect 52668 16210 52836 16212
rect 52668 16158 52670 16210
rect 52722 16158 52836 16210
rect 52668 16156 52836 16158
rect 52668 16146 52724 16156
rect 49756 16100 49812 16110
rect 49644 16098 49812 16100
rect 49644 16046 49758 16098
rect 49810 16046 49812 16098
rect 49644 16044 49812 16046
rect 46956 13748 47012 14588
rect 47964 15708 48356 15764
rect 49196 15874 49252 15886
rect 49196 15822 49198 15874
rect 49250 15822 49252 15874
rect 47516 14532 47572 14542
rect 47964 14532 48020 15708
rect 48412 15428 48468 15438
rect 48188 15426 48468 15428
rect 48188 15374 48414 15426
rect 48466 15374 48468 15426
rect 48188 15372 48468 15374
rect 48188 14642 48244 15372
rect 48412 15362 48468 15372
rect 49196 15428 49252 15822
rect 49196 15362 49252 15372
rect 49644 15316 49700 16044
rect 49756 16034 49812 16044
rect 50540 15988 50596 15998
rect 50540 15894 50596 15932
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50316 15428 50372 15438
rect 50316 15334 50372 15372
rect 49644 15314 50260 15316
rect 49644 15262 49646 15314
rect 49698 15262 50260 15314
rect 49644 15260 50260 15262
rect 49644 15250 49700 15260
rect 50204 15204 50260 15260
rect 52444 15204 52500 15214
rect 50204 15148 50820 15204
rect 48188 14590 48190 14642
rect 48242 14590 48244 14642
rect 48188 14578 48244 14590
rect 50316 14644 50372 14654
rect 50316 14550 50372 14588
rect 50764 14642 50820 15148
rect 52444 15202 52724 15204
rect 52444 15150 52446 15202
rect 52498 15150 52724 15202
rect 52444 15148 52724 15150
rect 52444 15138 52500 15148
rect 52668 15090 52724 15148
rect 52668 15038 52670 15090
rect 52722 15038 52724 15090
rect 52668 15026 52724 15038
rect 50764 14590 50766 14642
rect 50818 14590 50820 14642
rect 50764 14578 50820 14590
rect 47516 14530 48020 14532
rect 47516 14478 47518 14530
rect 47570 14478 48020 14530
rect 47516 14476 48020 14478
rect 47516 14466 47572 14476
rect 46956 13616 47012 13692
rect 47852 13748 47908 13758
rect 47628 13076 47684 13086
rect 47628 12290 47684 13020
rect 47628 12238 47630 12290
rect 47682 12238 47684 12290
rect 47628 12226 47684 12238
rect 46844 11342 46846 11394
rect 46898 11342 46900 11394
rect 46844 11330 46900 11342
rect 47516 11396 47572 11406
rect 47516 11302 47572 11340
rect 46396 11284 46452 11294
rect 46396 11190 46452 11228
rect 47404 11284 47460 11294
rect 47404 11190 47460 11228
rect 40012 10782 40014 10834
rect 40066 10782 40068 10834
rect 40012 10770 40068 10782
rect 45948 11172 46004 11182
rect 39452 10724 39508 10734
rect 39452 10722 39620 10724
rect 39452 10670 39454 10722
rect 39506 10670 39620 10722
rect 39452 10668 39620 10670
rect 39452 10658 39508 10668
rect 39340 10612 39396 10622
rect 39228 10610 39396 10612
rect 39228 10558 39342 10610
rect 39394 10558 39396 10610
rect 39228 10556 39396 10558
rect 31948 9874 32004 9884
rect 32620 9938 32676 10108
rect 38332 10098 38388 10108
rect 38444 10386 38500 10398
rect 38780 10388 38836 10398
rect 38444 10334 38446 10386
rect 38498 10334 38500 10386
rect 32620 9886 32622 9938
rect 32674 9886 32676 9938
rect 32620 9874 32676 9886
rect 33068 9940 33124 9950
rect 33068 9846 33124 9884
rect 38332 9940 38388 9950
rect 38444 9940 38500 10334
rect 38332 9938 38500 9940
rect 38332 9886 38334 9938
rect 38386 9886 38500 9938
rect 38332 9884 38500 9886
rect 38668 10386 38836 10388
rect 38668 10334 38782 10386
rect 38834 10334 38836 10386
rect 38668 10332 38836 10334
rect 38332 9874 38388 9884
rect 29820 9774 29822 9826
rect 29874 9774 29876 9826
rect 27468 9102 27470 9154
rect 27522 9102 27524 9154
rect 27468 9090 27524 9102
rect 27132 8990 27134 9042
rect 27186 8990 27188 9042
rect 27132 8428 27188 8990
rect 27692 8428 27748 9772
rect 27804 9762 27860 9772
rect 25452 8372 25620 8428
rect 24780 8318 24782 8370
rect 24834 8318 24836 8370
rect 24780 8306 24836 8318
rect 24444 8194 24500 8204
rect 24668 7588 24724 7598
rect 24668 7494 24724 7532
rect 23660 7362 24052 7364
rect 23660 7310 23662 7362
rect 23714 7310 24052 7362
rect 23660 7308 24052 7310
rect 24556 7362 24612 7374
rect 24556 7310 24558 7362
rect 24610 7310 24612 7362
rect 23660 6132 23716 7308
rect 24444 7252 24500 7262
rect 24444 7158 24500 7196
rect 24556 6916 24612 7310
rect 25564 7362 25620 8372
rect 26908 8372 27188 8428
rect 27468 8372 27748 8428
rect 27804 9154 27860 9166
rect 27804 9102 27806 9154
rect 27858 9102 27860 9154
rect 27804 8482 27860 9102
rect 27804 8430 27806 8482
rect 27858 8430 27860 8482
rect 26908 8370 26964 8372
rect 26908 8318 26910 8370
rect 26962 8318 26964 8370
rect 26908 8306 26964 8318
rect 27468 8034 27524 8372
rect 27468 7982 27470 8034
rect 27522 7982 27524 8034
rect 26236 7588 26292 7598
rect 25564 7310 25566 7362
rect 25618 7310 25620 7362
rect 25564 7252 25620 7310
rect 25564 7186 25620 7196
rect 26012 7532 26236 7588
rect 23884 6860 24612 6916
rect 23884 6802 23940 6860
rect 23884 6750 23886 6802
rect 23938 6750 23940 6802
rect 23884 6738 23940 6750
rect 26012 6802 26068 7532
rect 26236 7494 26292 7532
rect 26572 7476 26628 7514
rect 26572 7410 26628 7420
rect 27132 7476 27188 7486
rect 27132 7362 27188 7420
rect 27132 7310 27134 7362
rect 27186 7310 27188 7362
rect 27132 7298 27188 7310
rect 26012 6750 26014 6802
rect 26066 6750 26068 6802
rect 26012 6738 26068 6750
rect 26572 7250 26628 7262
rect 26572 7198 26574 7250
rect 26626 7198 26628 7250
rect 26572 6692 26628 7198
rect 26796 7252 26852 7262
rect 26796 6802 26852 7196
rect 26796 6750 26798 6802
rect 26850 6750 26852 6802
rect 26796 6738 26852 6750
rect 27356 7252 27412 7262
rect 27356 6804 27412 7196
rect 27468 6916 27524 7982
rect 27804 7588 27860 8430
rect 27804 7522 27860 7532
rect 27916 8930 27972 8942
rect 27916 8878 27918 8930
rect 27970 8878 27972 8930
rect 27916 8372 27972 8878
rect 29820 8428 29876 9774
rect 37660 9826 37716 9838
rect 37660 9774 37662 9826
rect 37714 9774 37716 9826
rect 30492 9716 30548 9726
rect 30492 9714 30772 9716
rect 30492 9662 30494 9714
rect 30546 9662 30772 9714
rect 30492 9660 30772 9662
rect 30492 9650 30548 9660
rect 30716 9266 30772 9660
rect 30716 9214 30718 9266
rect 30770 9214 30772 9266
rect 30716 9202 30772 9214
rect 37660 9044 37716 9774
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 28028 8372 28084 8382
rect 29820 8372 29988 8428
rect 27916 8370 28084 8372
rect 27916 8318 28030 8370
rect 28082 8318 28084 8370
rect 27916 8316 28084 8318
rect 27916 7476 27972 8316
rect 28028 8306 28084 8316
rect 27916 7410 27972 7420
rect 29932 7700 29988 8372
rect 29932 7474 29988 7644
rect 30492 7700 30548 7710
rect 30492 7606 30548 7644
rect 29932 7422 29934 7474
rect 29986 7422 29988 7474
rect 29932 7410 29988 7422
rect 27804 7364 27860 7374
rect 27692 6916 27748 6926
rect 27468 6914 27748 6916
rect 27468 6862 27694 6914
rect 27746 6862 27748 6914
rect 27468 6860 27748 6862
rect 27692 6850 27748 6860
rect 27356 6748 27524 6804
rect 26572 6626 26628 6636
rect 27244 6692 27300 6702
rect 27244 6598 27300 6636
rect 27468 6690 27524 6748
rect 27468 6638 27470 6690
rect 27522 6638 27524 6690
rect 27468 6626 27524 6638
rect 27804 6690 27860 7308
rect 29260 7364 29316 7374
rect 29260 7270 29316 7308
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 27804 6638 27806 6690
rect 27858 6638 27860 6690
rect 27804 6626 27860 6638
rect 37660 6690 37716 8988
rect 38668 8930 38724 10332
rect 38780 10322 38836 10332
rect 38668 8878 38670 8930
rect 38722 8878 38724 8930
rect 38668 8866 38724 8878
rect 38780 10164 38836 10174
rect 38780 8034 38836 10108
rect 39228 8930 39284 10556
rect 39340 10546 39396 10556
rect 39452 10388 39508 10398
rect 39228 8878 39230 8930
rect 39282 8878 39284 8930
rect 39228 8866 39284 8878
rect 39340 10386 39508 10388
rect 39340 10334 39454 10386
rect 39506 10334 39508 10386
rect 39340 10332 39508 10334
rect 38780 7982 38782 8034
rect 38834 7982 38836 8034
rect 38220 7476 38276 7486
rect 38220 7382 38276 7420
rect 38780 7476 38836 7982
rect 38780 7410 38836 7420
rect 39228 7476 39284 7486
rect 38332 7362 38388 7374
rect 38332 7310 38334 7362
rect 38386 7310 38388 7362
rect 38332 6802 38388 7310
rect 38556 7364 38612 7374
rect 38556 7270 38612 7308
rect 39116 7364 39172 7374
rect 39116 7270 39172 7308
rect 38332 6750 38334 6802
rect 38386 6750 38388 6802
rect 38332 6738 38388 6750
rect 37660 6638 37662 6690
rect 37714 6638 37716 6690
rect 37660 6626 37716 6638
rect 23660 6066 23716 6076
rect 26236 6132 26292 6142
rect 26236 6038 26292 6076
rect 19852 6020 19908 6030
rect 19628 6018 19908 6020
rect 19628 5966 19854 6018
rect 19906 5966 19908 6018
rect 19628 5964 19908 5966
rect 19852 5954 19908 5964
rect 39228 6020 39284 7420
rect 39340 7474 39396 10332
rect 39452 10322 39508 10332
rect 39564 9940 39620 10668
rect 41804 10722 41860 10734
rect 42812 10724 42868 10734
rect 41804 10670 41806 10722
rect 41858 10670 41860 10722
rect 39452 9044 39508 9054
rect 39564 9044 39620 9884
rect 40460 9940 40516 9950
rect 40460 9846 40516 9884
rect 41804 9938 41860 10670
rect 41804 9886 41806 9938
rect 41858 9886 41860 9938
rect 41804 9874 41860 9886
rect 42588 10722 42868 10724
rect 42588 10670 42814 10722
rect 42866 10670 42868 10722
rect 42588 10668 42868 10670
rect 41020 9826 41076 9838
rect 41020 9774 41022 9826
rect 41074 9774 41076 9826
rect 39452 9042 39620 9044
rect 39452 8990 39454 9042
rect 39506 8990 39620 9042
rect 39452 8988 39620 8990
rect 40236 9044 40292 9054
rect 39452 8978 39508 8988
rect 40236 8950 40292 8988
rect 40684 9044 40740 9054
rect 40684 8950 40740 8988
rect 41020 9044 41076 9774
rect 42588 9154 42644 10668
rect 42812 10658 42868 10668
rect 45948 10722 46004 11116
rect 47180 11172 47236 11182
rect 47180 11078 47236 11116
rect 45948 10670 45950 10722
rect 46002 10670 46004 10722
rect 45948 10658 46004 10670
rect 46620 10722 46676 10734
rect 46620 10670 46622 10722
rect 46674 10670 46676 10722
rect 45164 10612 45220 10622
rect 43932 10610 45220 10612
rect 43932 10558 45166 10610
rect 45218 10558 45220 10610
rect 43932 10556 45220 10558
rect 43932 9938 43988 10556
rect 45164 10546 45220 10556
rect 43932 9886 43934 9938
rect 43986 9886 43988 9938
rect 43932 9874 43988 9886
rect 44716 10388 44772 10398
rect 42588 9102 42590 9154
rect 42642 9102 42644 9154
rect 42588 9090 42644 9102
rect 44380 9602 44436 9614
rect 44380 9550 44382 9602
rect 44434 9550 44436 9602
rect 41020 8978 41076 8988
rect 41804 9044 41860 9054
rect 41860 8988 41972 9044
rect 41804 8950 41860 8988
rect 39340 7422 39342 7474
rect 39394 7422 39396 7474
rect 39340 7410 39396 7422
rect 39788 7474 39844 7486
rect 39788 7422 39790 7474
rect 39842 7422 39844 7474
rect 39788 6692 39844 7422
rect 41916 7364 41972 8988
rect 44380 8932 44436 9550
rect 44380 8866 44436 8876
rect 44604 9268 44660 9278
rect 44604 8258 44660 9212
rect 44716 8930 44772 10332
rect 45388 10388 45444 10398
rect 45388 10294 45444 10332
rect 45612 10386 45668 10398
rect 45836 10388 45892 10398
rect 45612 10334 45614 10386
rect 45666 10334 45668 10386
rect 45612 10164 45668 10334
rect 45388 10108 45668 10164
rect 45724 10386 45892 10388
rect 45724 10334 45838 10386
rect 45890 10334 45892 10386
rect 45724 10332 45892 10334
rect 45164 10052 45220 10062
rect 45164 9268 45220 9996
rect 45164 9136 45220 9212
rect 44716 8878 44718 8930
rect 44770 8878 44772 8930
rect 44716 8866 44772 8878
rect 44604 8206 44606 8258
rect 44658 8206 44660 8258
rect 44604 8194 44660 8206
rect 42476 8146 42532 8158
rect 42476 8094 42478 8146
rect 42530 8094 42532 8146
rect 42476 7474 42532 8094
rect 43260 7588 43316 7598
rect 43260 7494 43316 7532
rect 42476 7422 42478 7474
rect 42530 7422 42532 7474
rect 42476 7364 42532 7422
rect 41916 7362 42532 7364
rect 41916 7310 41918 7362
rect 41970 7310 42532 7362
rect 41916 7308 42532 7310
rect 45388 7362 45444 10108
rect 45500 9940 45556 9950
rect 45724 9940 45780 10332
rect 45836 10322 45892 10332
rect 45500 9938 45780 9940
rect 45500 9886 45502 9938
rect 45554 9886 45780 9938
rect 45500 9884 45780 9886
rect 46620 9940 46676 10670
rect 47852 10052 47908 13692
rect 47964 12180 48020 14476
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 52780 13748 52836 16156
rect 52892 15540 52948 17388
rect 53452 15988 53508 15998
rect 53452 15894 53508 15932
rect 53340 15540 53396 15550
rect 53676 15540 53732 18622
rect 54796 18562 54852 18574
rect 54796 18510 54798 18562
rect 54850 18510 54852 18562
rect 53788 18226 53844 18238
rect 53788 18174 53790 18226
rect 53842 18174 53844 18226
rect 53788 17778 53844 18174
rect 53788 17726 53790 17778
rect 53842 17726 53844 17778
rect 53788 17714 53844 17726
rect 54796 17780 54852 18510
rect 54796 17714 54852 17724
rect 55916 17780 55972 17790
rect 55916 17686 55972 17724
rect 56812 17780 56868 19180
rect 57148 17780 57204 17790
rect 56812 17778 57204 17780
rect 56812 17726 57150 17778
rect 57202 17726 57204 17778
rect 56812 17724 57204 17726
rect 56700 17668 56756 17678
rect 56812 17668 56868 17724
rect 57148 17714 57204 17724
rect 56700 17666 56868 17668
rect 56700 17614 56702 17666
rect 56754 17614 56868 17666
rect 56700 17612 56868 17614
rect 56700 17602 56756 17612
rect 52892 15538 53396 15540
rect 52892 15486 52894 15538
rect 52946 15486 53342 15538
rect 53394 15486 53396 15538
rect 52892 15484 53396 15486
rect 52892 15474 52948 15484
rect 53340 15474 53396 15484
rect 53452 15484 53732 15540
rect 53452 15316 53508 15484
rect 53228 15260 53508 15316
rect 54124 15426 54180 15438
rect 54124 15374 54126 15426
rect 54178 15374 54180 15426
rect 52780 13682 52836 13692
rect 53116 14644 53172 14654
rect 53116 13746 53172 14588
rect 53116 13694 53118 13746
rect 53170 13694 53172 13746
rect 53116 13682 53172 13694
rect 48412 13074 48468 13086
rect 48412 13022 48414 13074
rect 48466 13022 48468 13074
rect 48412 12404 48468 13022
rect 53228 12964 53284 15260
rect 53340 15090 53396 15102
rect 53340 15038 53342 15090
rect 53394 15038 53396 15090
rect 53340 13746 53396 15038
rect 53452 14644 53508 14654
rect 54124 14644 54180 15374
rect 53452 14642 53844 14644
rect 53452 14590 53454 14642
rect 53506 14590 53844 14642
rect 53452 14588 53844 14590
rect 53452 14578 53508 14588
rect 53676 13970 53732 13982
rect 53676 13918 53678 13970
rect 53730 13918 53732 13970
rect 53340 13694 53342 13746
rect 53394 13694 53396 13746
rect 53340 13682 53396 13694
rect 53564 13748 53620 13758
rect 53564 13654 53620 13692
rect 53452 12964 53508 12974
rect 53228 12962 53508 12964
rect 53228 12910 53454 12962
rect 53506 12910 53508 12962
rect 53228 12908 53508 12910
rect 53452 12898 53508 12908
rect 53676 12962 53732 13918
rect 53788 13746 53844 14588
rect 54124 14578 54180 14588
rect 55580 14644 55636 14654
rect 55580 14550 55636 14588
rect 53788 13694 53790 13746
rect 53842 13694 53844 13746
rect 53788 13682 53844 13694
rect 56364 14532 56420 14542
rect 56812 14532 56868 14542
rect 56364 14530 56868 14532
rect 56364 14478 56366 14530
rect 56418 14478 56814 14530
rect 56866 14478 56868 14530
rect 56364 14476 56868 14478
rect 53676 12910 53678 12962
rect 53730 12910 53732 12962
rect 53676 12898 53732 12910
rect 54124 12850 54180 12862
rect 54124 12798 54126 12850
rect 54178 12798 54180 12850
rect 48412 12338 48468 12348
rect 48860 12738 48916 12750
rect 48860 12686 48862 12738
rect 48914 12686 48916 12738
rect 48412 12180 48468 12190
rect 48860 12180 48916 12686
rect 52220 12740 52276 12750
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 49532 12292 49588 12302
rect 47964 12178 48916 12180
rect 47964 12126 48414 12178
rect 48466 12126 48916 12178
rect 47964 12124 48916 12126
rect 48972 12290 49588 12292
rect 48972 12238 49534 12290
rect 49586 12238 49588 12290
rect 48972 12236 49588 12238
rect 48412 12114 48468 12124
rect 48860 11508 48916 11518
rect 48972 11508 49028 12236
rect 49532 12226 49588 12236
rect 50764 12066 50820 12078
rect 50764 12014 50766 12066
rect 50818 12014 50820 12066
rect 50764 11620 50820 12014
rect 50764 11554 50820 11564
rect 51996 11732 52052 11742
rect 48860 11506 49028 11508
rect 48860 11454 48862 11506
rect 48914 11454 49028 11506
rect 48860 11452 49028 11454
rect 50988 11508 51044 11518
rect 48860 11442 48916 11452
rect 50988 11414 51044 11452
rect 48188 11394 48244 11406
rect 48188 11342 48190 11394
rect 48242 11342 48244 11394
rect 47852 9986 47908 9996
rect 48076 10052 48132 10062
rect 45500 9874 45556 9884
rect 46620 9874 46676 9884
rect 47628 9940 47684 9950
rect 47628 9846 47684 9884
rect 48076 9266 48132 9996
rect 48188 9828 48244 11342
rect 51996 11396 52052 11676
rect 51996 11302 52052 11340
rect 52220 11282 52276 12684
rect 53340 12740 53396 12750
rect 53340 12646 53396 12684
rect 53900 12740 53956 12750
rect 53900 12738 54068 12740
rect 53900 12686 53902 12738
rect 53954 12686 54068 12738
rect 53900 12684 54068 12686
rect 53900 12674 53956 12684
rect 53676 12404 53732 12414
rect 53676 12178 53732 12348
rect 53676 12126 53678 12178
rect 53730 12126 53732 12178
rect 53676 12114 53732 12126
rect 52892 12068 52948 12078
rect 52332 12066 52948 12068
rect 52332 12014 52894 12066
rect 52946 12014 52948 12066
rect 52332 12012 52948 12014
rect 52332 11618 52388 12012
rect 52892 12002 52948 12012
rect 52332 11566 52334 11618
rect 52386 11566 52388 11618
rect 52332 11554 52388 11566
rect 53564 11620 53620 11630
rect 53564 11526 53620 11564
rect 53676 11508 53732 11518
rect 53676 11414 53732 11452
rect 52220 11230 52222 11282
rect 52274 11230 52276 11282
rect 52220 11218 52276 11230
rect 53452 11396 53508 11406
rect 51436 11172 51492 11182
rect 51436 11170 51604 11172
rect 51436 11118 51438 11170
rect 51490 11118 51604 11170
rect 51436 11116 51604 11118
rect 51436 11106 51492 11116
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 48636 10722 48692 10734
rect 48636 10670 48638 10722
rect 48690 10670 48692 10722
rect 48300 9828 48356 9838
rect 48188 9826 48356 9828
rect 48188 9774 48302 9826
rect 48354 9774 48356 9826
rect 48188 9772 48356 9774
rect 48300 9380 48356 9772
rect 48636 9604 48692 10670
rect 50876 10612 50932 10622
rect 50876 10498 50932 10556
rect 51436 10612 51492 10622
rect 51436 10518 51492 10556
rect 50876 10446 50878 10498
rect 50930 10446 50932 10498
rect 50876 10052 50932 10446
rect 49532 9826 49588 9838
rect 49532 9774 49534 9826
rect 49586 9774 49588 9826
rect 48636 9538 48692 9548
rect 48860 9604 48916 9614
rect 49532 9604 49588 9774
rect 48860 9602 49588 9604
rect 48860 9550 48862 9602
rect 48914 9550 49588 9602
rect 48860 9548 49588 9550
rect 50316 9714 50372 9726
rect 50316 9662 50318 9714
rect 50370 9662 50372 9714
rect 50316 9604 50372 9662
rect 48860 9380 48916 9548
rect 48300 9324 48916 9380
rect 48076 9214 48078 9266
rect 48130 9214 48132 9266
rect 48076 9202 48132 9214
rect 48748 9154 48804 9166
rect 48748 9102 48750 9154
rect 48802 9102 48804 9154
rect 48748 8260 48804 9102
rect 48748 8194 48804 8204
rect 48972 8428 49028 9548
rect 50316 9538 50372 9548
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50876 9042 50932 9996
rect 50876 8990 50878 9042
rect 50930 8990 50932 9042
rect 50876 8978 50932 8990
rect 51548 8930 51604 11116
rect 52444 10164 52500 10174
rect 52444 9938 52500 10108
rect 52444 9886 52446 9938
rect 52498 9886 52500 9938
rect 52444 9874 52500 9886
rect 53452 9938 53508 11340
rect 53900 11394 53956 11406
rect 53900 11342 53902 11394
rect 53954 11342 53956 11394
rect 53900 10164 53956 11342
rect 53900 10098 53956 10108
rect 53452 9886 53454 9938
rect 53506 9886 53508 9938
rect 53452 9874 53508 9886
rect 51548 8878 51550 8930
rect 51602 8878 51604 8930
rect 51548 8428 51604 8878
rect 48972 8372 49140 8428
rect 48972 8258 49028 8372
rect 49084 8306 49140 8316
rect 51324 8372 51604 8428
rect 54012 8428 54068 12684
rect 54124 11620 54180 12798
rect 54460 12740 54516 12750
rect 54460 12402 54516 12684
rect 54460 12350 54462 12402
rect 54514 12350 54516 12402
rect 54460 12338 54516 12350
rect 55020 12404 55076 12414
rect 55020 12310 55076 12348
rect 56364 12404 56420 14476
rect 56812 14466 56868 14476
rect 54236 11954 54292 11966
rect 54236 11902 54238 11954
rect 54290 11902 54292 11954
rect 54236 11844 54292 11902
rect 54236 11778 54292 11788
rect 54572 11954 54628 11966
rect 54572 11902 54574 11954
rect 54626 11902 54628 11954
rect 54236 11620 54292 11630
rect 54124 11618 54292 11620
rect 54124 11566 54238 11618
rect 54290 11566 54292 11618
rect 54124 11564 54292 11566
rect 54236 11554 54292 11564
rect 54124 11396 54180 11406
rect 54124 11302 54180 11340
rect 51772 8372 51828 8382
rect 51324 8306 51380 8316
rect 48972 8206 48974 8258
rect 49026 8206 49028 8258
rect 45500 8034 45556 8046
rect 47180 8036 47236 8046
rect 45500 7982 45502 8034
rect 45554 7982 45556 8034
rect 45500 7588 45556 7982
rect 45500 7522 45556 7532
rect 46956 8034 47236 8036
rect 46956 7982 47182 8034
rect 47234 7982 47236 8034
rect 46956 7980 47236 7982
rect 45388 7310 45390 7362
rect 45442 7310 45444 7362
rect 40460 6802 40516 6814
rect 40460 6750 40462 6802
rect 40514 6750 40516 6802
rect 39788 6626 39844 6636
rect 40012 6692 40068 6702
rect 40012 6130 40068 6636
rect 40460 6692 40516 6750
rect 40460 6626 40516 6636
rect 40012 6078 40014 6130
rect 40066 6078 40068 6130
rect 40012 6066 40068 6078
rect 40908 6466 40964 6478
rect 40908 6414 40910 6466
rect 40962 6414 40964 6466
rect 39788 6020 39844 6030
rect 39228 6018 39844 6020
rect 39228 5966 39230 6018
rect 39282 5966 39790 6018
rect 39842 5966 39844 6018
rect 39228 5964 39844 5966
rect 39228 5954 39284 5964
rect 39788 5954 39844 5964
rect 19180 5854 19182 5906
rect 19234 5854 19236 5906
rect 19180 5842 19236 5854
rect 1820 5794 1876 5806
rect 1820 5742 1822 5794
rect 1874 5742 1876 5794
rect 28 3668 84 3678
rect 28 800 84 3612
rect 1820 3554 1876 5742
rect 21980 5794 22036 5806
rect 21980 5742 21982 5794
rect 22034 5742 22036 5794
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 2492 3668 2548 3678
rect 2492 3574 2548 3612
rect 21532 3668 21588 3678
rect 1820 3502 1822 3554
rect 1874 3502 1876 3554
rect 1820 3490 1876 3502
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 21532 800 21588 3612
rect 21980 3554 22036 5742
rect 40124 5682 40180 5694
rect 40124 5630 40126 5682
rect 40178 5630 40180 5682
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 40124 5236 40180 5630
rect 40124 5170 40180 5180
rect 40572 5124 40628 5134
rect 40572 5030 40628 5068
rect 40908 5124 40964 6414
rect 41244 5236 41300 5246
rect 41244 5142 41300 5180
rect 40908 5058 40964 5068
rect 41916 5124 41972 7308
rect 45388 7298 45444 7310
rect 46284 6804 46340 6814
rect 46284 6690 46340 6748
rect 46284 6638 46286 6690
rect 46338 6638 46340 6690
rect 46284 6626 46340 6638
rect 46956 6690 47012 7980
rect 47180 7970 47236 7980
rect 48972 6804 49028 8206
rect 49756 8260 49812 8270
rect 49756 8166 49812 8204
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 51772 7698 51828 8316
rect 51884 8370 51940 8382
rect 51884 8318 51886 8370
rect 51938 8318 51940 8370
rect 51884 8260 51940 8318
rect 51884 8194 51940 8204
rect 52668 8372 52724 8382
rect 54012 8372 54404 8428
rect 51772 7646 51774 7698
rect 51826 7646 51828 7698
rect 51772 7634 51828 7646
rect 50428 7586 50484 7598
rect 50428 7534 50430 7586
rect 50482 7534 50484 7586
rect 48972 6738 49028 6748
rect 49084 6802 49140 6814
rect 49084 6750 49086 6802
rect 49138 6750 49140 6802
rect 46956 6638 46958 6690
rect 47010 6638 47012 6690
rect 46956 6626 47012 6638
rect 49084 6692 49140 6750
rect 49084 6626 49140 6636
rect 49420 6804 49476 6814
rect 49420 6130 49476 6748
rect 49644 6804 49700 6814
rect 49644 6690 49700 6748
rect 50428 6802 50484 7534
rect 52332 7364 52388 7374
rect 52332 7270 52388 7308
rect 50428 6750 50430 6802
rect 50482 6750 50484 6802
rect 50428 6738 50484 6750
rect 52556 6916 52612 6926
rect 52556 6802 52612 6860
rect 52556 6750 52558 6802
rect 52610 6750 52612 6802
rect 52556 6738 52612 6750
rect 52668 6804 52724 8316
rect 53564 8258 53620 8270
rect 53564 8206 53566 8258
rect 53618 8206 53620 8258
rect 53564 7364 53620 8206
rect 53564 7298 53620 7308
rect 53788 8258 53844 8270
rect 53788 8206 53790 8258
rect 53842 8206 53844 8258
rect 53788 6916 53844 8206
rect 53788 6850 53844 6860
rect 54012 8258 54068 8270
rect 54012 8206 54014 8258
rect 54066 8206 54068 8258
rect 49644 6638 49646 6690
rect 49698 6638 49700 6690
rect 49644 6626 49700 6638
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 49420 6078 49422 6130
rect 49474 6078 49476 6130
rect 49420 6066 49476 6078
rect 52668 6132 52724 6748
rect 53340 6804 53396 6814
rect 52780 6132 52836 6142
rect 52668 6130 52836 6132
rect 52668 6078 52782 6130
rect 52834 6078 52836 6130
rect 52668 6076 52836 6078
rect 52780 6066 52836 6076
rect 53340 5906 53396 6748
rect 54012 6692 54068 8206
rect 54124 8260 54180 8270
rect 54124 8166 54180 8204
rect 54124 8036 54180 8046
rect 54348 8036 54404 8372
rect 54124 8034 54404 8036
rect 54124 7982 54126 8034
rect 54178 7982 54404 8034
rect 54124 7980 54404 7982
rect 54124 7970 54180 7980
rect 54460 7588 54516 7598
rect 54460 7494 54516 7532
rect 54572 7140 54628 11902
rect 54908 11170 54964 11182
rect 54908 11118 54910 11170
rect 54962 11118 54964 11170
rect 54908 9940 54964 11118
rect 56364 10722 56420 12348
rect 56364 10670 56366 10722
rect 56418 10670 56420 10722
rect 54908 9874 54964 9884
rect 55580 9940 55636 9950
rect 55580 9846 55636 9884
rect 56364 9940 56420 10670
rect 56812 9940 56868 9950
rect 56364 9938 56868 9940
rect 56364 9886 56814 9938
rect 56866 9886 56868 9938
rect 56364 9884 56868 9886
rect 56364 9826 56420 9884
rect 56812 9874 56868 9884
rect 56364 9774 56366 9826
rect 56418 9774 56420 9826
rect 55356 9154 55412 9166
rect 55356 9102 55358 9154
rect 55410 9102 55412 9154
rect 55244 7700 55300 7710
rect 55244 7474 55300 7644
rect 55356 7588 55412 9102
rect 56364 8428 56420 9774
rect 56252 8372 56420 8428
rect 55692 7700 55748 7710
rect 55692 7606 55748 7644
rect 56252 7700 56308 8372
rect 56252 7634 56308 7644
rect 55356 7522 55412 7532
rect 55244 7422 55246 7474
rect 55298 7422 55300 7474
rect 55244 7410 55300 7422
rect 54012 6626 54068 6636
rect 54124 7084 54628 7140
rect 54124 6018 54180 7084
rect 54124 5966 54126 6018
rect 54178 5966 54180 6018
rect 54124 5954 54180 5966
rect 53340 5854 53342 5906
rect 53394 5854 53396 5906
rect 53340 5842 53396 5854
rect 56252 5794 56308 5806
rect 56252 5742 56254 5794
rect 56306 5742 56308 5794
rect 55356 5460 55412 5470
rect 41916 5058 41972 5068
rect 43372 5234 43428 5246
rect 43372 5182 43374 5234
rect 43426 5182 43428 5234
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 22428 3668 22484 3678
rect 22428 3574 22484 3612
rect 21980 3502 21982 3554
rect 22034 3502 22036 3554
rect 21980 3490 22036 3502
rect 43372 3556 43428 5182
rect 55356 5234 55412 5404
rect 55356 5182 55358 5234
rect 55410 5182 55412 5234
rect 55356 5170 55412 5182
rect 43932 5124 43988 5134
rect 43932 5030 43988 5068
rect 56140 5124 56196 5134
rect 56252 5124 56308 5742
rect 56140 5122 56308 5124
rect 56140 5070 56142 5122
rect 56194 5070 56308 5122
rect 56140 5068 56308 5070
rect 56140 5058 56196 5068
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 43372 3490 43428 3500
rect 43708 3668 43764 3678
rect 43708 800 43764 3612
rect 45612 3668 45668 3678
rect 45612 3574 45668 3612
rect 44940 3556 44996 3566
rect 44940 3462 44996 3500
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 0 200 112 800
rect 21504 200 21616 800
rect 43680 200 43792 800
<< via2 >>
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4172 51884 4228 51940
rect 2044 50706 2100 50708
rect 2044 50654 2046 50706
rect 2046 50654 2098 50706
rect 2098 50654 2100 50706
rect 2044 50652 2100 50654
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4284 50540 4340 50596
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 8316 52162 8372 52164
rect 8316 52110 8318 52162
rect 8318 52110 8370 52162
rect 8370 52110 8372 52162
rect 8316 52108 8372 52110
rect 8876 52108 8932 52164
rect 8428 51938 8484 51940
rect 8428 51886 8430 51938
rect 8430 51886 8482 51938
rect 8482 51886 8484 51938
rect 8428 51884 8484 51886
rect 8540 51772 8596 51828
rect 5068 50652 5124 50708
rect 4956 50594 5012 50596
rect 4956 50542 4958 50594
rect 4958 50542 5010 50594
rect 5010 50542 5012 50594
rect 4956 50540 5012 50542
rect 6524 50594 6580 50596
rect 6524 50542 6526 50594
rect 6526 50542 6578 50594
rect 6578 50542 6580 50594
rect 6524 50540 6580 50542
rect 7308 49980 7364 50036
rect 8764 49868 8820 49924
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 7308 49026 7364 49028
rect 7308 48974 7310 49026
rect 7310 48974 7362 49026
rect 7362 48974 7364 49026
rect 7308 48972 7364 48974
rect 7532 48636 7588 48692
rect 4956 48300 5012 48356
rect 7308 48354 7364 48356
rect 7308 48302 7310 48354
rect 7310 48302 7362 48354
rect 7362 48302 7364 48354
rect 7308 48300 7364 48302
rect 7420 48242 7476 48244
rect 7420 48190 7422 48242
rect 7422 48190 7474 48242
rect 7474 48190 7476 48242
rect 7420 48188 7476 48190
rect 7980 48748 8036 48804
rect 8316 48636 8372 48692
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 7868 47570 7924 47572
rect 7868 47518 7870 47570
rect 7870 47518 7922 47570
rect 7922 47518 7924 47570
rect 7868 47516 7924 47518
rect 7644 47180 7700 47236
rect 7308 47068 7364 47124
rect 2828 46002 2884 46004
rect 2828 45950 2830 46002
rect 2830 45950 2882 46002
rect 2882 45950 2884 46002
rect 2828 45948 2884 45950
rect 5740 46786 5796 46788
rect 5740 46734 5742 46786
rect 5742 46734 5794 46786
rect 5794 46734 5796 46786
rect 5740 46732 5796 46734
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 3500 45948 3556 46004
rect 4956 46002 5012 46004
rect 4956 45950 4958 46002
rect 4958 45950 5010 46002
rect 5010 45950 5012 46002
rect 4956 45948 5012 45950
rect 8540 48972 8596 49028
rect 8652 48802 8708 48804
rect 8652 48750 8654 48802
rect 8654 48750 8706 48802
rect 8706 48750 8708 48802
rect 8652 48748 8708 48750
rect 8764 48636 8820 48692
rect 9100 52162 9156 52164
rect 9100 52110 9102 52162
rect 9102 52110 9154 52162
rect 9154 52110 9156 52162
rect 9100 52108 9156 52110
rect 9324 51772 9380 51828
rect 8988 51378 9044 51380
rect 8988 51326 8990 51378
rect 8990 51326 9042 51378
rect 9042 51326 9044 51378
rect 8988 51324 9044 51326
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 9772 51378 9828 51380
rect 9772 51326 9774 51378
rect 9774 51326 9826 51378
rect 9826 51326 9828 51378
rect 9772 51324 9828 51326
rect 14140 51324 14196 51380
rect 10108 50594 10164 50596
rect 10108 50542 10110 50594
rect 10110 50542 10162 50594
rect 10162 50542 10164 50594
rect 10108 50540 10164 50542
rect 12012 50540 12068 50596
rect 9884 50034 9940 50036
rect 9884 49982 9886 50034
rect 9886 49982 9938 50034
rect 9938 49982 9940 50034
rect 9884 49980 9940 49982
rect 10780 49980 10836 50036
rect 11676 50034 11732 50036
rect 11676 49982 11678 50034
rect 11678 49982 11730 50034
rect 11730 49982 11732 50034
rect 11676 49980 11732 49982
rect 9772 49922 9828 49924
rect 9772 49870 9774 49922
rect 9774 49870 9826 49922
rect 9826 49870 9828 49922
rect 9772 49868 9828 49870
rect 8428 47180 8484 47236
rect 8316 47068 8372 47124
rect 8652 47516 8708 47572
rect 8988 48188 9044 48244
rect 11900 49810 11956 49812
rect 11900 49758 11902 49810
rect 11902 49758 11954 49810
rect 11954 49758 11956 49810
rect 11900 49756 11956 49758
rect 10108 49532 10164 49588
rect 9660 48242 9716 48244
rect 9660 48190 9662 48242
rect 9662 48190 9714 48242
rect 9714 48190 9716 48242
rect 9660 48188 9716 48190
rect 11564 49586 11620 49588
rect 11564 49534 11566 49586
rect 11566 49534 11618 49586
rect 11618 49534 11620 49586
rect 11564 49532 11620 49534
rect 10780 48076 10836 48132
rect 8764 47180 8820 47236
rect 8652 46956 8708 47012
rect 8988 46786 9044 46788
rect 8988 46734 8990 46786
rect 8990 46734 9042 46786
rect 9042 46734 9044 46786
rect 8988 46732 9044 46734
rect 5068 45612 5124 45668
rect 5404 45948 5460 46004
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4172 43708 4228 43764
rect 2156 41916 2212 41972
rect 3052 30882 3108 30884
rect 3052 30830 3054 30882
rect 3054 30830 3106 30882
rect 3106 30830 3108 30882
rect 3052 30828 3108 30830
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4396 41970 4452 41972
rect 4396 41918 4398 41970
rect 4398 41918 4450 41970
rect 4450 41918 4452 41970
rect 4396 41916 4452 41918
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5628 45666 5684 45668
rect 5628 45614 5630 45666
rect 5630 45614 5682 45666
rect 5682 45614 5684 45666
rect 5628 45612 5684 45614
rect 5852 45612 5908 45668
rect 8092 45666 8148 45668
rect 8092 45614 8094 45666
rect 8094 45614 8146 45666
rect 8146 45614 8148 45666
rect 8092 45612 8148 45614
rect 10220 47180 10276 47236
rect 9884 46674 9940 46676
rect 9884 46622 9886 46674
rect 9886 46622 9938 46674
rect 9938 46622 9940 46674
rect 9884 46620 9940 46622
rect 11900 47234 11956 47236
rect 11900 47182 11902 47234
rect 11902 47182 11954 47234
rect 11954 47182 11956 47234
rect 11900 47180 11956 47182
rect 12460 49980 12516 50036
rect 13244 50540 13300 50596
rect 13692 49980 13748 50036
rect 13916 50428 13972 50484
rect 12684 49756 12740 49812
rect 13580 49586 13636 49588
rect 13580 49534 13582 49586
rect 13582 49534 13634 49586
rect 13634 49534 13636 49586
rect 13580 49532 13636 49534
rect 12460 48188 12516 48244
rect 12908 48802 12964 48804
rect 12908 48750 12910 48802
rect 12910 48750 12962 48802
rect 12962 48750 12964 48802
rect 12908 48748 12964 48750
rect 13132 48748 13188 48804
rect 12796 48242 12852 48244
rect 12796 48190 12798 48242
rect 12798 48190 12850 48242
rect 12850 48190 12852 48242
rect 12796 48188 12852 48190
rect 13804 48748 13860 48804
rect 14028 48748 14084 48804
rect 13244 48188 13300 48244
rect 12908 48130 12964 48132
rect 12908 48078 12910 48130
rect 12910 48078 12962 48130
rect 12962 48078 12964 48130
rect 12908 48076 12964 48078
rect 12012 46620 12068 46676
rect 12908 46620 12964 46676
rect 13692 46508 13748 46564
rect 13580 46002 13636 46004
rect 13580 45950 13582 46002
rect 13582 45950 13634 46002
rect 13634 45950 13636 46002
rect 13580 45948 13636 45950
rect 12908 45836 12964 45892
rect 9884 45052 9940 45108
rect 5852 44268 5908 44324
rect 6412 44322 6468 44324
rect 6412 44270 6414 44322
rect 6414 44270 6466 44322
rect 6466 44270 6468 44322
rect 6412 44268 6468 44270
rect 9996 44268 10052 44324
rect 10444 45106 10500 45108
rect 10444 45054 10446 45106
rect 10446 45054 10498 45106
rect 10498 45054 10500 45106
rect 10444 45052 10500 45054
rect 13916 48242 13972 48244
rect 13916 48190 13918 48242
rect 13918 48190 13970 48242
rect 13970 48190 13972 48242
rect 13916 48188 13972 48190
rect 14364 50540 14420 50596
rect 15820 50482 15876 50484
rect 15820 50430 15822 50482
rect 15822 50430 15874 50482
rect 15874 50430 15876 50482
rect 15820 50428 15876 50430
rect 16604 50428 16660 50484
rect 17052 50482 17108 50484
rect 17052 50430 17054 50482
rect 17054 50430 17106 50482
rect 17106 50430 17108 50482
rect 17052 50428 17108 50430
rect 17948 50428 18004 50484
rect 17276 48972 17332 49028
rect 18508 50428 18564 50484
rect 19628 50428 19684 50484
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19964 49868 20020 49924
rect 20972 49868 21028 49924
rect 20748 49138 20804 49140
rect 20748 49086 20750 49138
rect 20750 49086 20802 49138
rect 20802 49086 20804 49138
rect 20748 49084 20804 49086
rect 14140 46732 14196 46788
rect 14140 45948 14196 46004
rect 13916 45836 13972 45892
rect 10332 44322 10388 44324
rect 10332 44270 10334 44322
rect 10334 44270 10386 44322
rect 10386 44270 10388 44322
rect 10332 44268 10388 44270
rect 9324 43484 9380 43540
rect 8316 43372 8372 43428
rect 6188 43260 6244 43316
rect 5852 41916 5908 41972
rect 5068 41804 5124 41860
rect 5628 41858 5684 41860
rect 5628 41806 5630 41858
rect 5630 41806 5682 41858
rect 5682 41806 5684 41858
rect 5628 41804 5684 41806
rect 6076 41916 6132 41972
rect 9884 43314 9940 43316
rect 9884 43262 9886 43314
rect 9886 43262 9938 43314
rect 9938 43262 9940 43314
rect 9884 43260 9940 43262
rect 16828 46844 16884 46900
rect 15036 46732 15092 46788
rect 14476 45890 14532 45892
rect 14476 45838 14478 45890
rect 14478 45838 14530 45890
rect 14530 45838 14532 45890
rect 14476 45836 14532 45838
rect 10220 43538 10276 43540
rect 10220 43486 10222 43538
rect 10222 43486 10274 43538
rect 10274 43486 10276 43538
rect 10220 43484 10276 43486
rect 10108 42924 10164 42980
rect 8428 41916 8484 41972
rect 9324 41916 9380 41972
rect 9996 41916 10052 41972
rect 10332 41916 10388 41972
rect 10780 43426 10836 43428
rect 10780 43374 10782 43426
rect 10782 43374 10834 43426
rect 10834 43374 10836 43426
rect 10780 43372 10836 43374
rect 15372 46562 15428 46564
rect 15372 46510 15374 46562
rect 15374 46510 15426 46562
rect 15426 46510 15428 46562
rect 15372 46508 15428 46510
rect 17612 46898 17668 46900
rect 17612 46846 17614 46898
rect 17614 46846 17666 46898
rect 17666 46846 17668 46898
rect 17612 46844 17668 46846
rect 16940 46786 16996 46788
rect 16940 46734 16942 46786
rect 16942 46734 16994 46786
rect 16994 46734 16996 46786
rect 16940 46732 16996 46734
rect 17388 46060 17444 46116
rect 16828 45836 16884 45892
rect 17164 45836 17220 45892
rect 16380 45388 16436 45444
rect 15260 45276 15316 45332
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 24444 50428 24500 50484
rect 21980 49868 22036 49924
rect 24892 49868 24948 49924
rect 24220 49532 24276 49588
rect 21868 49138 21924 49140
rect 21868 49086 21870 49138
rect 21870 49086 21922 49138
rect 21922 49086 21924 49138
rect 21868 49084 21924 49086
rect 22988 49138 23044 49140
rect 22988 49086 22990 49138
rect 22990 49086 23042 49138
rect 23042 49086 23044 49138
rect 22988 49084 23044 49086
rect 21644 49026 21700 49028
rect 21644 48974 21646 49026
rect 21646 48974 21698 49026
rect 21698 48974 21700 49026
rect 21644 48972 21700 48974
rect 21644 47682 21700 47684
rect 21644 47630 21646 47682
rect 21646 47630 21698 47682
rect 21698 47630 21700 47682
rect 21644 47628 21700 47630
rect 23212 48300 23268 48356
rect 23212 47628 23268 47684
rect 18396 46732 18452 46788
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 18060 45388 18116 45444
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 17724 45330 17780 45332
rect 17724 45278 17726 45330
rect 17726 45278 17778 45330
rect 17778 45278 17780 45330
rect 17724 45276 17780 45278
rect 15036 43372 15092 43428
rect 14252 42978 14308 42980
rect 14252 42926 14254 42978
rect 14254 42926 14306 42978
rect 14306 42926 14308 42978
rect 14252 42924 14308 42926
rect 14588 42978 14644 42980
rect 14588 42926 14590 42978
rect 14590 42926 14642 42978
rect 14642 42926 14644 42978
rect 14588 42924 14644 42926
rect 12908 42866 12964 42868
rect 12908 42814 12910 42866
rect 12910 42814 12962 42866
rect 12962 42814 12964 42866
rect 12908 42812 12964 42814
rect 14812 42754 14868 42756
rect 14812 42702 14814 42754
rect 14814 42702 14866 42754
rect 14866 42702 14868 42754
rect 14812 42700 14868 42702
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 11676 41916 11732 41972
rect 10780 41020 10836 41076
rect 7756 38780 7812 38836
rect 9772 38834 9828 38836
rect 9772 38782 9774 38834
rect 9774 38782 9826 38834
rect 9826 38782 9828 38834
rect 9772 38780 9828 38782
rect 8316 38050 8372 38052
rect 8316 37998 8318 38050
rect 8318 37998 8370 38050
rect 8370 37998 8372 38050
rect 8316 37996 8372 37998
rect 7868 37436 7924 37492
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4508 35698 4564 35700
rect 4508 35646 4510 35698
rect 4510 35646 4562 35698
rect 4562 35646 4564 35698
rect 4508 35644 4564 35646
rect 7756 36706 7812 36708
rect 7756 36654 7758 36706
rect 7758 36654 7810 36706
rect 7810 36654 7812 36706
rect 7756 36652 7812 36654
rect 5404 35644 5460 35700
rect 8316 36652 8372 36708
rect 8764 37490 8820 37492
rect 8764 37438 8766 37490
rect 8766 37438 8818 37490
rect 8818 37438 8820 37490
rect 8764 37436 8820 37438
rect 13580 41916 13636 41972
rect 15036 41970 15092 41972
rect 15036 41918 15038 41970
rect 15038 41918 15090 41970
rect 15090 41918 15092 41970
rect 15036 41916 15092 41918
rect 11676 41132 11732 41188
rect 12348 41186 12404 41188
rect 12348 41134 12350 41186
rect 12350 41134 12402 41186
rect 12402 41134 12404 41186
rect 12348 41132 12404 41134
rect 11788 41074 11844 41076
rect 11788 41022 11790 41074
rect 11790 41022 11842 41074
rect 11842 41022 11844 41074
rect 11788 41020 11844 41022
rect 13020 40514 13076 40516
rect 13020 40462 13022 40514
rect 13022 40462 13074 40514
rect 13074 40462 13076 40514
rect 13020 40460 13076 40462
rect 13692 40460 13748 40516
rect 15036 40348 15092 40404
rect 10892 37436 10948 37492
rect 11228 37490 11284 37492
rect 11228 37438 11230 37490
rect 11230 37438 11282 37490
rect 11282 37438 11284 37490
rect 11228 37436 11284 37438
rect 11788 37436 11844 37492
rect 12684 38162 12740 38164
rect 12684 38110 12686 38162
rect 12686 38110 12738 38162
rect 12738 38110 12740 38162
rect 12684 38108 12740 38110
rect 13356 38108 13412 38164
rect 7980 36594 8036 36596
rect 7980 36542 7982 36594
rect 7982 36542 8034 36594
rect 8034 36542 8036 36594
rect 7980 36540 8036 36542
rect 9100 36594 9156 36596
rect 9100 36542 9102 36594
rect 9102 36542 9154 36594
rect 9154 36542 9156 36594
rect 9100 36540 9156 36542
rect 7756 35698 7812 35700
rect 7756 35646 7758 35698
rect 7758 35646 7810 35698
rect 7810 35646 7812 35698
rect 7756 35644 7812 35646
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 12460 35644 12516 35700
rect 13244 35698 13300 35700
rect 13244 35646 13246 35698
rect 13246 35646 13298 35698
rect 13298 35646 13300 35698
rect 13244 35644 13300 35646
rect 20188 45388 20244 45444
rect 23436 48188 23492 48244
rect 24780 49586 24836 49588
rect 24780 49534 24782 49586
rect 24782 49534 24834 49586
rect 24834 49534 24836 49586
rect 24780 49532 24836 49534
rect 25900 50428 25956 50484
rect 25788 49922 25844 49924
rect 25788 49870 25790 49922
rect 25790 49870 25842 49922
rect 25842 49870 25844 49922
rect 25788 49868 25844 49870
rect 25116 49644 25172 49700
rect 25676 49698 25732 49700
rect 25676 49646 25678 49698
rect 25678 49646 25730 49698
rect 25730 49646 25732 49698
rect 25676 49644 25732 49646
rect 24892 49084 24948 49140
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 26236 50428 26292 50484
rect 27692 50428 27748 50484
rect 26460 49698 26516 49700
rect 26460 49646 26462 49698
rect 26462 49646 26514 49698
rect 26514 49646 26516 49698
rect 26460 49644 26516 49646
rect 25116 48914 25172 48916
rect 25116 48862 25118 48914
rect 25118 48862 25170 48914
rect 25170 48862 25172 48914
rect 25116 48860 25172 48862
rect 24668 48466 24724 48468
rect 24668 48414 24670 48466
rect 24670 48414 24722 48466
rect 24722 48414 24724 48466
rect 24668 48412 24724 48414
rect 24444 48354 24500 48356
rect 24444 48302 24446 48354
rect 24446 48302 24498 48354
rect 24498 48302 24500 48354
rect 24444 48300 24500 48302
rect 24332 48242 24388 48244
rect 24332 48190 24334 48242
rect 24334 48190 24386 48242
rect 24386 48190 24388 48242
rect 24332 48188 24388 48190
rect 24332 47570 24388 47572
rect 24332 47518 24334 47570
rect 24334 47518 24386 47570
rect 24386 47518 24388 47570
rect 24332 47516 24388 47518
rect 25564 48412 25620 48468
rect 21756 46114 21812 46116
rect 21756 46062 21758 46114
rect 21758 46062 21810 46114
rect 21810 46062 21812 46114
rect 21756 46060 21812 46062
rect 20860 46002 20916 46004
rect 20860 45950 20862 46002
rect 20862 45950 20914 46002
rect 20914 45950 20916 46002
rect 20860 45948 20916 45950
rect 21868 46002 21924 46004
rect 21868 45950 21870 46002
rect 21870 45950 21922 46002
rect 21922 45950 21924 46002
rect 21868 45948 21924 45950
rect 21644 45388 21700 45444
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 18060 43484 18116 43540
rect 18396 43538 18452 43540
rect 18396 43486 18398 43538
rect 18398 43486 18450 43538
rect 18450 43486 18452 43538
rect 18396 43484 18452 43486
rect 16044 42924 16100 42980
rect 15484 42812 15540 42868
rect 15596 42700 15652 42756
rect 15036 38108 15092 38164
rect 14700 37996 14756 38052
rect 15484 38050 15540 38052
rect 15484 37998 15486 38050
rect 15486 37998 15538 38050
rect 15538 37998 15540 38050
rect 15484 37996 15540 37998
rect 18844 43484 18900 43540
rect 20188 43484 20244 43540
rect 20860 44322 20916 44324
rect 20860 44270 20862 44322
rect 20862 44270 20914 44322
rect 20914 44270 20916 44322
rect 20860 44268 20916 44270
rect 16492 42194 16548 42196
rect 16492 42142 16494 42194
rect 16494 42142 16546 42194
rect 16546 42142 16548 42194
rect 16492 42140 16548 42142
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 17500 42140 17556 42196
rect 21756 44322 21812 44324
rect 21756 44270 21758 44322
rect 21758 44270 21810 44322
rect 21810 44270 21812 44322
rect 21756 44268 21812 44270
rect 21196 43426 21252 43428
rect 21196 43374 21198 43426
rect 21198 43374 21250 43426
rect 21250 43374 21252 43426
rect 21196 43372 21252 43374
rect 23212 45388 23268 45444
rect 22540 44210 22596 44212
rect 22540 44158 22542 44210
rect 22542 44158 22594 44210
rect 22594 44158 22596 44210
rect 22540 44156 22596 44158
rect 22092 43372 22148 43428
rect 23548 42866 23604 42868
rect 23548 42814 23550 42866
rect 23550 42814 23602 42866
rect 23602 42814 23604 42866
rect 23548 42812 23604 42814
rect 15820 41970 15876 41972
rect 15820 41918 15822 41970
rect 15822 41918 15874 41970
rect 15874 41918 15876 41970
rect 15820 41916 15876 41918
rect 19404 41970 19460 41972
rect 19404 41918 19406 41970
rect 19406 41918 19458 41970
rect 19458 41918 19460 41970
rect 19404 41916 19460 41918
rect 17164 41132 17220 41188
rect 17724 41186 17780 41188
rect 17724 41134 17726 41186
rect 17726 41134 17778 41186
rect 17778 41134 17780 41186
rect 17724 41132 17780 41134
rect 19404 41132 19460 41188
rect 20300 41916 20356 41972
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19964 40460 20020 40516
rect 19068 40402 19124 40404
rect 19068 40350 19070 40402
rect 19070 40350 19122 40402
rect 19122 40350 19124 40402
rect 19068 40348 19124 40350
rect 20860 41916 20916 41972
rect 20636 41298 20692 41300
rect 20636 41246 20638 41298
rect 20638 41246 20690 41298
rect 20690 41246 20692 41298
rect 20636 41244 20692 41246
rect 21868 41298 21924 41300
rect 21868 41246 21870 41298
rect 21870 41246 21922 41298
rect 21922 41246 21924 41298
rect 21868 41244 21924 41246
rect 21644 40460 21700 40516
rect 21084 40402 21140 40404
rect 21084 40350 21086 40402
rect 21086 40350 21138 40402
rect 21138 40350 21140 40402
rect 21084 40348 21140 40350
rect 22316 39618 22372 39620
rect 22316 39566 22318 39618
rect 22318 39566 22370 39618
rect 22370 39566 22372 39618
rect 22316 39564 22372 39566
rect 20300 39340 20356 39396
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 21532 39394 21588 39396
rect 21532 39342 21534 39394
rect 21534 39342 21586 39394
rect 21586 39342 21588 39394
rect 21532 39340 21588 39342
rect 24780 46562 24836 46564
rect 24780 46510 24782 46562
rect 24782 46510 24834 46562
rect 24834 46510 24836 46562
rect 24780 46508 24836 46510
rect 26684 49532 26740 49588
rect 26012 48412 26068 48468
rect 25676 48130 25732 48132
rect 25676 48078 25678 48130
rect 25678 48078 25730 48130
rect 25730 48078 25732 48130
rect 25676 48076 25732 48078
rect 26572 48914 26628 48916
rect 26572 48862 26574 48914
rect 26574 48862 26626 48914
rect 26626 48862 26628 48914
rect 26572 48860 26628 48862
rect 27356 49644 27412 49700
rect 27020 48636 27076 48692
rect 26348 48076 26404 48132
rect 25676 47516 25732 47572
rect 24668 45836 24724 45892
rect 24108 45276 24164 45332
rect 24668 44828 24724 44884
rect 26908 46620 26964 46676
rect 26124 46562 26180 46564
rect 26124 46510 26126 46562
rect 26126 46510 26178 46562
rect 26178 46510 26180 46562
rect 26124 46508 26180 46510
rect 25564 45164 25620 45220
rect 26796 45890 26852 45892
rect 26796 45838 26798 45890
rect 26798 45838 26850 45890
rect 26850 45838 26852 45890
rect 26796 45836 26852 45838
rect 25788 44828 25844 44884
rect 25900 45052 25956 45108
rect 24892 44492 24948 44548
rect 25452 44546 25508 44548
rect 25452 44494 25454 44546
rect 25454 44494 25506 44546
rect 25506 44494 25508 44546
rect 25452 44492 25508 44494
rect 26236 45106 26292 45108
rect 26236 45054 26238 45106
rect 26238 45054 26290 45106
rect 26290 45054 26292 45106
rect 26236 45052 26292 45054
rect 26012 44716 26068 44772
rect 26124 44492 26180 44548
rect 26684 45330 26740 45332
rect 26684 45278 26686 45330
rect 26686 45278 26738 45330
rect 26738 45278 26740 45330
rect 26684 45276 26740 45278
rect 26908 44604 26964 44660
rect 27244 44546 27300 44548
rect 27244 44494 27246 44546
rect 27246 44494 27298 44546
rect 27298 44494 27300 44546
rect 27244 44492 27300 44494
rect 26796 44210 26852 44212
rect 26796 44158 26798 44210
rect 26798 44158 26850 44210
rect 26850 44158 26852 44210
rect 26796 44156 26852 44158
rect 25788 42194 25844 42196
rect 25788 42142 25790 42194
rect 25790 42142 25842 42194
rect 25842 42142 25844 42194
rect 25788 42140 25844 42142
rect 26124 42812 26180 42868
rect 26572 42194 26628 42196
rect 26572 42142 26574 42194
rect 26574 42142 26626 42194
rect 26626 42142 26628 42194
rect 26572 42140 26628 42142
rect 26460 41916 26516 41972
rect 23212 41074 23268 41076
rect 23212 41022 23214 41074
rect 23214 41022 23266 41074
rect 23266 41022 23268 41074
rect 23212 41020 23268 41022
rect 22988 40460 23044 40516
rect 22764 39340 22820 39396
rect 14476 35644 14532 35700
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 16156 36540 16212 36596
rect 17388 36594 17444 36596
rect 17388 36542 17390 36594
rect 17390 36542 17442 36594
rect 17442 36542 17444 36594
rect 17388 36540 17444 36542
rect 16604 35698 16660 35700
rect 16604 35646 16606 35698
rect 16606 35646 16658 35698
rect 16658 35646 16660 35698
rect 16604 35644 16660 35646
rect 17612 35698 17668 35700
rect 17612 35646 17614 35698
rect 17614 35646 17666 35698
rect 17666 35646 17668 35698
rect 17612 35644 17668 35646
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 17948 35644 18004 35700
rect 18284 35644 18340 35700
rect 13692 34860 13748 34916
rect 8204 34748 8260 34804
rect 8988 34748 9044 34804
rect 6188 33964 6244 34020
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 5964 31052 6020 31108
rect 14252 34914 14308 34916
rect 14252 34862 14254 34914
rect 14254 34862 14306 34914
rect 14306 34862 14308 34914
rect 14252 34860 14308 34862
rect 15036 34860 15092 34916
rect 9772 34018 9828 34020
rect 9772 33966 9774 34018
rect 9774 33966 9826 34018
rect 9826 33966 9828 34018
rect 9772 33964 9828 33966
rect 12236 33964 12292 34020
rect 6188 31052 6244 31108
rect 6412 31106 6468 31108
rect 6412 31054 6414 31106
rect 6414 31054 6466 31106
rect 6466 31054 6468 31106
rect 6412 31052 6468 31054
rect 10108 31106 10164 31108
rect 10108 31054 10110 31106
rect 10110 31054 10162 31106
rect 10162 31054 10164 31106
rect 10108 31052 10164 31054
rect 5068 30828 5124 30884
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 28700 4228 28756
rect 5180 28588 5236 28644
rect 5404 28476 5460 28532
rect 5964 28476 6020 28532
rect 6188 28642 6244 28644
rect 6188 28590 6190 28642
rect 6190 28590 6242 28642
rect 6242 28590 6244 28642
rect 6188 28588 6244 28590
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 2716 23436 2772 23492
rect 4172 26178 4228 26180
rect 4172 26126 4174 26178
rect 4174 26126 4226 26178
rect 4226 26126 4228 26178
rect 4172 26124 4228 26126
rect 6188 26124 6244 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 8988 29426 9044 29428
rect 8988 29374 8990 29426
rect 8990 29374 9042 29426
rect 9042 29374 9044 29426
rect 8988 29372 9044 29374
rect 9660 29372 9716 29428
rect 6636 28812 6692 28868
rect 7532 28866 7588 28868
rect 7532 28814 7534 28866
rect 7534 28814 7586 28866
rect 7586 28814 7588 28866
rect 7532 28812 7588 28814
rect 8204 28812 8260 28868
rect 7308 28530 7364 28532
rect 7308 28478 7310 28530
rect 7310 28478 7362 28530
rect 7362 28478 7364 28530
rect 7308 28476 7364 28478
rect 6524 26796 6580 26852
rect 6300 25730 6356 25732
rect 6300 25678 6302 25730
rect 6302 25678 6354 25730
rect 6354 25678 6356 25730
rect 6300 25676 6356 25678
rect 6860 26850 6916 26852
rect 6860 26798 6862 26850
rect 6862 26798 6914 26850
rect 6914 26798 6916 26850
rect 6860 26796 6916 26798
rect 7532 26796 7588 26852
rect 7308 26348 7364 26404
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 3388 23436 3444 23492
rect 3948 23436 4004 23492
rect 2268 21868 2324 21924
rect 6076 23212 6132 23268
rect 6972 25676 7028 25732
rect 12908 32732 12964 32788
rect 13804 32732 13860 32788
rect 14364 31836 14420 31892
rect 12908 31164 12964 31220
rect 16492 34188 16548 34244
rect 15484 34076 15540 34132
rect 15036 30994 15092 30996
rect 15036 30942 15038 30994
rect 15038 30942 15090 30994
rect 15090 30942 15092 30994
rect 15036 30940 15092 30942
rect 15372 30940 15428 30996
rect 12236 29596 12292 29652
rect 13132 29650 13188 29652
rect 13132 29598 13134 29650
rect 13134 29598 13186 29650
rect 13186 29598 13188 29650
rect 13132 29596 13188 29598
rect 9436 28364 9492 28420
rect 16716 34130 16772 34132
rect 16716 34078 16718 34130
rect 16718 34078 16770 34130
rect 16770 34078 16772 34130
rect 16716 34076 16772 34078
rect 17724 34242 17780 34244
rect 17724 34190 17726 34242
rect 17726 34190 17778 34242
rect 17778 34190 17780 34242
rect 17724 34188 17780 34190
rect 21196 35698 21252 35700
rect 21196 35646 21198 35698
rect 21198 35646 21250 35698
rect 21250 35646 21252 35698
rect 21196 35644 21252 35646
rect 22988 35532 23044 35588
rect 20860 35084 20916 35140
rect 22428 35138 22484 35140
rect 22428 35086 22430 35138
rect 22430 35086 22482 35138
rect 22482 35086 22484 35138
rect 22428 35084 22484 35086
rect 26908 41020 26964 41076
rect 24332 40460 24388 40516
rect 23548 39340 23604 39396
rect 24556 39564 24612 39620
rect 26684 40402 26740 40404
rect 26684 40350 26686 40402
rect 26686 40350 26738 40402
rect 26738 40350 26740 40402
rect 26684 40348 26740 40350
rect 25676 39730 25732 39732
rect 25676 39678 25678 39730
rect 25678 39678 25730 39730
rect 25730 39678 25732 39730
rect 25676 39676 25732 39678
rect 25564 39564 25620 39620
rect 25116 38780 25172 38836
rect 24220 37490 24276 37492
rect 24220 37438 24222 37490
rect 24222 37438 24274 37490
rect 24274 37438 24276 37490
rect 24220 37436 24276 37438
rect 27468 46674 27524 46676
rect 27468 46622 27470 46674
rect 27470 46622 27522 46674
rect 27522 46622 27524 46674
rect 27468 46620 27524 46622
rect 33964 50428 34020 50484
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 28700 48914 28756 48916
rect 28700 48862 28702 48914
rect 28702 48862 28754 48914
rect 28754 48862 28756 48914
rect 28700 48860 28756 48862
rect 30044 48914 30100 48916
rect 30044 48862 30046 48914
rect 30046 48862 30098 48914
rect 30098 48862 30100 48914
rect 30044 48860 30100 48862
rect 27692 46620 27748 46676
rect 27804 48636 27860 48692
rect 27804 47292 27860 47348
rect 28476 47346 28532 47348
rect 28476 47294 28478 47346
rect 28478 47294 28530 47346
rect 28530 47294 28532 47346
rect 28476 47292 28532 47294
rect 28700 47404 28756 47460
rect 30268 47404 30324 47460
rect 30716 47458 30772 47460
rect 30716 47406 30718 47458
rect 30718 47406 30770 47458
rect 30770 47406 30772 47458
rect 30716 47404 30772 47406
rect 29484 47346 29540 47348
rect 29484 47294 29486 47346
rect 29486 47294 29538 47346
rect 29538 47294 29540 47346
rect 29484 47292 29540 47294
rect 33852 48802 33908 48804
rect 33852 48750 33854 48802
rect 33854 48750 33906 48802
rect 33906 48750 33908 48802
rect 33852 48748 33908 48750
rect 30940 47292 30996 47348
rect 29820 47180 29876 47236
rect 27916 45836 27972 45892
rect 28476 46674 28532 46676
rect 28476 46622 28478 46674
rect 28478 46622 28530 46674
rect 28530 46622 28532 46674
rect 28476 46620 28532 46622
rect 27916 45388 27972 45444
rect 28140 45388 28196 45444
rect 28476 45388 28532 45444
rect 29820 45666 29876 45668
rect 29820 45614 29822 45666
rect 29822 45614 29874 45666
rect 29874 45614 29876 45666
rect 29820 45612 29876 45614
rect 28812 45276 28868 45332
rect 28140 45106 28196 45108
rect 28140 45054 28142 45106
rect 28142 45054 28194 45106
rect 28194 45054 28196 45106
rect 28140 45052 28196 45054
rect 28364 44940 28420 44996
rect 29708 44940 29764 44996
rect 28924 44434 28980 44436
rect 28924 44382 28926 44434
rect 28926 44382 28978 44434
rect 28978 44382 28980 44434
rect 28924 44380 28980 44382
rect 30604 45500 30660 45556
rect 30268 45106 30324 45108
rect 30268 45054 30270 45106
rect 30270 45054 30322 45106
rect 30322 45054 30324 45106
rect 30268 45052 30324 45054
rect 30828 46002 30884 46004
rect 30828 45950 30830 46002
rect 30830 45950 30882 46002
rect 30882 45950 30884 46002
rect 30828 45948 30884 45950
rect 31276 46562 31332 46564
rect 31276 46510 31278 46562
rect 31278 46510 31330 46562
rect 31330 46510 31332 46562
rect 31276 46508 31332 46510
rect 31276 45948 31332 46004
rect 31164 45388 31220 45444
rect 29932 44434 29988 44436
rect 29932 44382 29934 44434
rect 29934 44382 29986 44434
rect 29986 44382 29988 44434
rect 29932 44380 29988 44382
rect 30156 44322 30212 44324
rect 30156 44270 30158 44322
rect 30158 44270 30210 44322
rect 30210 44270 30212 44322
rect 30156 44268 30212 44270
rect 30828 44322 30884 44324
rect 30828 44270 30830 44322
rect 30830 44270 30882 44322
rect 30882 44270 30884 44322
rect 30828 44268 30884 44270
rect 31388 45500 31444 45556
rect 32172 47458 32228 47460
rect 32172 47406 32174 47458
rect 32174 47406 32226 47458
rect 32226 47406 32228 47458
rect 32172 47404 32228 47406
rect 32508 47404 32564 47460
rect 31836 47346 31892 47348
rect 31836 47294 31838 47346
rect 31838 47294 31890 47346
rect 31890 47294 31892 47346
rect 31836 47292 31892 47294
rect 31948 47234 32004 47236
rect 31948 47182 31950 47234
rect 31950 47182 32002 47234
rect 32002 47182 32004 47234
rect 31948 47180 32004 47182
rect 36316 50428 36372 50484
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 36876 49810 36932 49812
rect 36876 49758 36878 49810
rect 36878 49758 36930 49810
rect 36930 49758 36932 49810
rect 36876 49756 36932 49758
rect 34412 48748 34468 48804
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 36540 47628 36596 47684
rect 36764 47570 36820 47572
rect 36764 47518 36766 47570
rect 36766 47518 36818 47570
rect 36818 47518 36820 47570
rect 36764 47516 36820 47518
rect 37436 50428 37492 50484
rect 39452 50482 39508 50484
rect 39452 50430 39454 50482
rect 39454 50430 39506 50482
rect 39506 50430 39508 50482
rect 39452 50428 39508 50430
rect 40012 50428 40068 50484
rect 40348 50428 40404 50484
rect 37660 50370 37716 50372
rect 37660 50318 37662 50370
rect 37662 50318 37714 50370
rect 37714 50318 37716 50370
rect 37660 50316 37716 50318
rect 39676 50316 39732 50372
rect 42252 49810 42308 49812
rect 42252 49758 42254 49810
rect 42254 49758 42306 49810
rect 42306 49758 42308 49810
rect 42252 49756 42308 49758
rect 37772 47682 37828 47684
rect 37772 47630 37774 47682
rect 37774 47630 37826 47682
rect 37826 47630 37828 47682
rect 37772 47628 37828 47630
rect 37996 47570 38052 47572
rect 37996 47518 37998 47570
rect 37998 47518 38050 47570
rect 38050 47518 38052 47570
rect 37996 47516 38052 47518
rect 40796 48130 40852 48132
rect 40796 48078 40798 48130
rect 40798 48078 40850 48130
rect 40850 48078 40852 48130
rect 40796 48076 40852 48078
rect 38332 46956 38388 47012
rect 41580 47068 41636 47124
rect 32732 46508 32788 46564
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 41692 46956 41748 47012
rect 32956 45612 33012 45668
rect 37660 45890 37716 45892
rect 37660 45838 37662 45890
rect 37662 45838 37714 45890
rect 37714 45838 37716 45890
rect 37660 45836 37716 45838
rect 31724 45388 31780 45444
rect 27804 42140 27860 42196
rect 40796 45836 40852 45892
rect 41020 45890 41076 45892
rect 41020 45838 41022 45890
rect 41022 45838 41074 45890
rect 41074 45838 41076 45890
rect 41020 45836 41076 45838
rect 41468 45836 41524 45892
rect 40796 45330 40852 45332
rect 40796 45278 40798 45330
rect 40798 45278 40850 45330
rect 40850 45278 40852 45330
rect 40796 45276 40852 45278
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 31612 42028 31668 42084
rect 29260 41970 29316 41972
rect 29260 41918 29262 41970
rect 29262 41918 29314 41970
rect 29314 41918 29316 41970
rect 29260 41916 29316 41918
rect 27244 40402 27300 40404
rect 27244 40350 27246 40402
rect 27246 40350 27298 40402
rect 27298 40350 27300 40402
rect 27244 40348 27300 40350
rect 28588 40460 28644 40516
rect 27020 39676 27076 39732
rect 26796 38834 26852 38836
rect 26796 38782 26798 38834
rect 26798 38782 26850 38834
rect 26850 38782 26852 38834
rect 26796 38780 26852 38782
rect 27692 39564 27748 39620
rect 32060 41356 32116 41412
rect 33628 42028 33684 42084
rect 29260 40514 29316 40516
rect 29260 40462 29262 40514
rect 29262 40462 29314 40514
rect 29314 40462 29316 40514
rect 29260 40460 29316 40462
rect 34748 42082 34804 42084
rect 34748 42030 34750 42082
rect 34750 42030 34802 42082
rect 34802 42030 34804 42082
rect 34748 42028 34804 42030
rect 34412 41298 34468 41300
rect 34412 41246 34414 41298
rect 34414 41246 34466 41298
rect 34466 41246 34468 41298
rect 34412 41244 34468 41246
rect 29708 39618 29764 39620
rect 29708 39566 29710 39618
rect 29710 39566 29762 39618
rect 29762 39566 29764 39618
rect 29708 39564 29764 39566
rect 27692 38780 27748 38836
rect 26684 37436 26740 37492
rect 24892 36540 24948 36596
rect 25340 36594 25396 36596
rect 25340 36542 25342 36594
rect 25342 36542 25394 36594
rect 25394 36542 25396 36594
rect 25340 36540 25396 36542
rect 28364 38834 28420 38836
rect 28364 38782 28366 38834
rect 28366 38782 28418 38834
rect 28418 38782 28420 38834
rect 28364 38780 28420 38782
rect 31612 38834 31668 38836
rect 31612 38782 31614 38834
rect 31614 38782 31666 38834
rect 31666 38782 31668 38834
rect 31612 38780 31668 38782
rect 32172 39564 32228 39620
rect 32956 39618 33012 39620
rect 32956 39566 32958 39618
rect 32958 39566 33010 39618
rect 33010 39566 33012 39618
rect 32956 39564 33012 39566
rect 32844 38892 32900 38948
rect 33628 38946 33684 38948
rect 33628 38894 33630 38946
rect 33630 38894 33682 38946
rect 33682 38894 33684 38946
rect 33628 38892 33684 38894
rect 40460 45052 40516 45108
rect 38108 44994 38164 44996
rect 38108 44942 38110 44994
rect 38110 44942 38162 44994
rect 38162 44942 38164 44994
rect 38108 44940 38164 44942
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35756 42028 35812 42084
rect 36988 42028 37044 42084
rect 36540 41970 36596 41972
rect 36540 41918 36542 41970
rect 36542 41918 36594 41970
rect 36594 41918 36596 41970
rect 36540 41916 36596 41918
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 41410 35252 41412
rect 35196 41358 35198 41410
rect 35198 41358 35250 41410
rect 35250 41358 35252 41410
rect 35196 41356 35252 41358
rect 35308 41298 35364 41300
rect 35308 41246 35310 41298
rect 35310 41246 35362 41298
rect 35362 41246 35364 41298
rect 35308 41244 35364 41246
rect 35644 40236 35700 40292
rect 40236 43484 40292 43540
rect 38108 42028 38164 42084
rect 38780 41916 38836 41972
rect 37884 40402 37940 40404
rect 37884 40350 37886 40402
rect 37886 40350 37938 40402
rect 37938 40350 37940 40402
rect 37884 40348 37940 40350
rect 39340 42028 39396 42084
rect 38780 40348 38836 40404
rect 37324 40236 37380 40292
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35084 38834 35140 38836
rect 35084 38782 35086 38834
rect 35086 38782 35138 38834
rect 35138 38782 35140 38834
rect 35084 38780 35140 38782
rect 36988 38722 37044 38724
rect 36988 38670 36990 38722
rect 36990 38670 37042 38722
rect 37042 38670 37044 38722
rect 36988 38668 37044 38670
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34972 38162 35028 38164
rect 34972 38110 34974 38162
rect 34974 38110 35026 38162
rect 35026 38110 35028 38162
rect 34972 38108 35028 38110
rect 36316 38162 36372 38164
rect 36316 38110 36318 38162
rect 36318 38110 36370 38162
rect 36370 38110 36372 38162
rect 36316 38108 36372 38110
rect 36652 38162 36708 38164
rect 36652 38110 36654 38162
rect 36654 38110 36706 38162
rect 36706 38110 36708 38162
rect 36652 38108 36708 38110
rect 34636 37378 34692 37380
rect 34636 37326 34638 37378
rect 34638 37326 34690 37378
rect 34690 37326 34692 37378
rect 34636 37324 34692 37326
rect 36764 37938 36820 37940
rect 36764 37886 36766 37938
rect 36766 37886 36818 37938
rect 36818 37886 36820 37938
rect 36764 37884 36820 37886
rect 35532 37324 35588 37380
rect 32172 37212 32228 37268
rect 33852 37266 33908 37268
rect 33852 37214 33854 37266
rect 33854 37214 33906 37266
rect 33906 37214 33908 37266
rect 33852 37212 33908 37214
rect 35084 37212 35140 37268
rect 32508 37154 32564 37156
rect 32508 37102 32510 37154
rect 32510 37102 32562 37154
rect 32562 37102 32564 37154
rect 32508 37100 32564 37102
rect 23548 35644 23604 35700
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 18732 34130 18788 34132
rect 18732 34078 18734 34130
rect 18734 34078 18786 34130
rect 18786 34078 18788 34130
rect 18732 34076 18788 34078
rect 16156 32786 16212 32788
rect 16156 32734 16158 32786
rect 16158 32734 16210 32786
rect 16210 32734 16212 32786
rect 16156 32732 16212 32734
rect 17164 32732 17220 32788
rect 15708 31836 15764 31892
rect 17948 31836 18004 31892
rect 16268 31164 16324 31220
rect 18508 30994 18564 30996
rect 18508 30942 18510 30994
rect 18510 30942 18562 30994
rect 18562 30942 18564 30994
rect 18508 30940 18564 30942
rect 15148 28418 15204 28420
rect 15148 28366 15150 28418
rect 15150 28366 15202 28418
rect 15202 28366 15204 28418
rect 15148 28364 15204 28366
rect 12908 27356 12964 27412
rect 7532 26124 7588 26180
rect 7980 26348 8036 26404
rect 7868 26066 7924 26068
rect 7868 26014 7870 26066
rect 7870 26014 7922 26066
rect 7922 26014 7924 26066
rect 7868 26012 7924 26014
rect 10108 26908 10164 26964
rect 11228 26908 11284 26964
rect 8764 26066 8820 26068
rect 8764 26014 8766 26066
rect 8766 26014 8818 26066
rect 8818 26014 8820 26066
rect 8764 26012 8820 26014
rect 9996 26402 10052 26404
rect 9996 26350 9998 26402
rect 9998 26350 10050 26402
rect 10050 26350 10052 26402
rect 9996 26348 10052 26350
rect 9772 26066 9828 26068
rect 9772 26014 9774 26066
rect 9774 26014 9826 26066
rect 9826 26014 9828 26066
rect 9772 26012 9828 26014
rect 8204 25676 8260 25732
rect 12908 27186 12964 27188
rect 12908 27134 12910 27186
rect 12910 27134 12962 27186
rect 12962 27134 12964 27186
rect 12908 27132 12964 27134
rect 14924 27692 14980 27748
rect 14700 27356 14756 27412
rect 14812 27186 14868 27188
rect 14812 27134 14814 27186
rect 14814 27134 14866 27186
rect 14866 27134 14868 27186
rect 14812 27132 14868 27134
rect 13020 26908 13076 26964
rect 13580 26962 13636 26964
rect 13580 26910 13582 26962
rect 13582 26910 13634 26962
rect 13634 26910 13636 26962
rect 13580 26908 13636 26910
rect 7084 23548 7140 23604
rect 6860 23212 6916 23268
rect 8428 23212 8484 23268
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 2716 21868 2772 21924
rect 4732 21868 4788 21924
rect 4956 21868 5012 21924
rect 5628 21868 5684 21924
rect 2492 21532 2548 21588
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 2828 20524 2884 20580
rect 3836 20578 3892 20580
rect 3836 20526 3838 20578
rect 3838 20526 3890 20578
rect 3890 20526 3892 20578
rect 3836 20524 3892 20526
rect 6636 22988 6692 23044
rect 6076 21868 6132 21924
rect 8428 22482 8484 22484
rect 8428 22430 8430 22482
rect 8430 22430 8482 22482
rect 8482 22430 8484 22482
rect 8428 22428 8484 22430
rect 8988 22428 9044 22484
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 5068 19404 5124 19460
rect 4956 19346 5012 19348
rect 4956 19294 4958 19346
rect 4958 19294 5010 19346
rect 5010 19294 5012 19346
rect 4956 19292 5012 19294
rect 9100 22316 9156 22372
rect 11228 23378 11284 23380
rect 11228 23326 11230 23378
rect 11230 23326 11282 23378
rect 11282 23326 11284 23378
rect 11228 23324 11284 23326
rect 9660 23266 9716 23268
rect 9660 23214 9662 23266
rect 9662 23214 9714 23266
rect 9714 23214 9716 23266
rect 9660 23212 9716 23214
rect 11228 22988 11284 23044
rect 11788 23324 11844 23380
rect 9436 21532 9492 21588
rect 9884 21586 9940 21588
rect 9884 21534 9886 21586
rect 9886 21534 9938 21586
rect 9938 21534 9940 21586
rect 9884 21532 9940 21534
rect 6300 19458 6356 19460
rect 6300 19406 6302 19458
rect 6302 19406 6354 19458
rect 6354 19406 6356 19458
rect 6300 19404 6356 19406
rect 6748 19458 6804 19460
rect 6748 19406 6750 19458
rect 6750 19406 6802 19458
rect 6802 19406 6804 19458
rect 6748 19404 6804 19406
rect 8540 19404 8596 19460
rect 6076 19346 6132 19348
rect 6076 19294 6078 19346
rect 6078 19294 6130 19346
rect 6130 19294 6132 19346
rect 6076 19292 6132 19294
rect 2156 18396 2212 18452
rect 7868 18450 7924 18452
rect 7868 18398 7870 18450
rect 7870 18398 7922 18450
rect 7922 18398 7924 18450
rect 7868 18396 7924 18398
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 8316 17666 8372 17668
rect 8316 17614 8318 17666
rect 8318 17614 8370 17666
rect 8370 17614 8372 17666
rect 8316 17612 8372 17614
rect 5068 16716 5124 16772
rect 5740 16716 5796 16772
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 7980 15036 8036 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 1932 12012 1988 12068
rect 6300 13634 6356 13636
rect 6300 13582 6302 13634
rect 6302 13582 6354 13634
rect 6354 13582 6356 13634
rect 6300 13580 6356 13582
rect 6860 13634 6916 13636
rect 6860 13582 6862 13634
rect 6862 13582 6914 13634
rect 6914 13582 6916 13634
rect 6860 13580 6916 13582
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4172 13020 4228 13076
rect 6972 13074 7028 13076
rect 6972 13022 6974 13074
rect 6974 13022 7026 13074
rect 7026 13022 7028 13074
rect 6972 13020 7028 13022
rect 6076 12962 6132 12964
rect 6076 12910 6078 12962
rect 6078 12910 6130 12962
rect 6130 12910 6132 12962
rect 6076 12908 6132 12910
rect 7308 12908 7364 12964
rect 4284 12684 4340 12740
rect 3500 12012 3556 12068
rect 3948 12066 4004 12068
rect 3948 12014 3950 12066
rect 3950 12014 4002 12066
rect 4002 12014 4004 12066
rect 3948 12012 4004 12014
rect 3164 10610 3220 10612
rect 3164 10558 3166 10610
rect 3166 10558 3218 10610
rect 3218 10558 3220 10610
rect 3164 10556 3220 10558
rect 2828 10444 2884 10500
rect 2156 7532 2212 7588
rect 5740 12738 5796 12740
rect 5740 12686 5742 12738
rect 5742 12686 5794 12738
rect 5794 12686 5796 12738
rect 5740 12684 5796 12686
rect 6636 12684 6692 12740
rect 6860 12796 6916 12852
rect 7196 12348 7252 12404
rect 5740 12012 5796 12068
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 6524 11282 6580 11284
rect 6524 11230 6526 11282
rect 6526 11230 6578 11282
rect 6578 11230 6580 11282
rect 6524 11228 6580 11230
rect 4396 10610 4452 10612
rect 4396 10558 4398 10610
rect 4398 10558 4450 10610
rect 4450 10558 4452 10610
rect 4396 10556 4452 10558
rect 6748 11228 6804 11284
rect 7756 12908 7812 12964
rect 8204 12796 8260 12852
rect 7756 12738 7812 12740
rect 7756 12686 7758 12738
rect 7758 12686 7810 12738
rect 7810 12686 7812 12738
rect 7756 12684 7812 12686
rect 8988 16882 9044 16884
rect 8988 16830 8990 16882
rect 8990 16830 9042 16882
rect 9042 16830 9044 16882
rect 8988 16828 9044 16830
rect 12012 23154 12068 23156
rect 12012 23102 12014 23154
rect 12014 23102 12066 23154
rect 12066 23102 12068 23154
rect 12012 23100 12068 23102
rect 13020 23996 13076 24052
rect 12908 23826 12964 23828
rect 12908 23774 12910 23826
rect 12910 23774 12962 23826
rect 12962 23774 12964 23826
rect 12908 23772 12964 23774
rect 13020 23324 13076 23380
rect 15036 27298 15092 27300
rect 15036 27246 15038 27298
rect 15038 27246 15090 27298
rect 15090 27246 15092 27298
rect 15036 27244 15092 27246
rect 14924 26908 14980 26964
rect 13356 23266 13412 23268
rect 13356 23214 13358 23266
rect 13358 23214 13410 23266
rect 13410 23214 13412 23266
rect 13356 23212 13412 23214
rect 12684 23154 12740 23156
rect 12684 23102 12686 23154
rect 12686 23102 12738 23154
rect 12738 23102 12740 23154
rect 12684 23100 12740 23102
rect 13132 23100 13188 23156
rect 12012 22370 12068 22372
rect 12012 22318 12014 22370
rect 12014 22318 12066 22370
rect 12066 22318 12068 22370
rect 12012 22316 12068 22318
rect 12348 20578 12404 20580
rect 12348 20526 12350 20578
rect 12350 20526 12402 20578
rect 12402 20526 12404 20578
rect 12348 20524 12404 20526
rect 14476 23826 14532 23828
rect 14476 23774 14478 23826
rect 14478 23774 14530 23826
rect 14530 23774 14532 23826
rect 14476 23772 14532 23774
rect 13804 23212 13860 23268
rect 14588 23324 14644 23380
rect 13580 23100 13636 23156
rect 14924 23324 14980 23380
rect 16380 30268 16436 30324
rect 16716 30268 16772 30324
rect 18620 30268 18676 30324
rect 19404 31890 19460 31892
rect 19404 31838 19406 31890
rect 19406 31838 19458 31890
rect 19458 31838 19460 31890
rect 19404 31836 19460 31838
rect 20748 33628 20804 33684
rect 22428 33628 22484 33684
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 24444 35698 24500 35700
rect 24444 35646 24446 35698
rect 24446 35646 24498 35698
rect 24498 35646 24500 35698
rect 24444 35644 24500 35646
rect 31500 36988 31556 37044
rect 27916 35644 27972 35700
rect 23996 35586 24052 35588
rect 23996 35534 23998 35586
rect 23998 35534 24050 35586
rect 24050 35534 24052 35586
rect 23996 35532 24052 35534
rect 19628 31836 19684 31892
rect 19292 31500 19348 31556
rect 19068 30994 19124 30996
rect 19068 30942 19070 30994
rect 19070 30942 19122 30994
rect 19122 30942 19124 30994
rect 19068 30940 19124 30942
rect 19180 30380 19236 30436
rect 20300 31554 20356 31556
rect 20300 31502 20302 31554
rect 20302 31502 20354 31554
rect 20354 31502 20356 31554
rect 20300 31500 20356 31502
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20188 30434 20244 30436
rect 20188 30382 20190 30434
rect 20190 30382 20242 30434
rect 20242 30382 20244 30434
rect 20188 30380 20244 30382
rect 20300 30268 20356 30324
rect 20076 30210 20132 30212
rect 20076 30158 20078 30210
rect 20078 30158 20130 30210
rect 20130 30158 20132 30210
rect 20076 30156 20132 30158
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 18732 28700 18788 28756
rect 19516 28476 19572 28532
rect 20860 31890 20916 31892
rect 20860 31838 20862 31890
rect 20862 31838 20914 31890
rect 20914 31838 20916 31890
rect 20860 31836 20916 31838
rect 24892 32450 24948 32452
rect 24892 32398 24894 32450
rect 24894 32398 24946 32450
rect 24946 32398 24948 32450
rect 24892 32396 24948 32398
rect 20524 30156 20580 30212
rect 20412 28476 20468 28532
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 15708 28028 15764 28084
rect 21644 30322 21700 30324
rect 21644 30270 21646 30322
rect 21646 30270 21698 30322
rect 21698 30270 21700 30322
rect 21644 30268 21700 30270
rect 28588 35698 28644 35700
rect 28588 35646 28590 35698
rect 28590 35646 28642 35698
rect 28642 35646 28644 35698
rect 28588 35644 28644 35646
rect 32172 37042 32228 37044
rect 32172 36990 32174 37042
rect 32174 36990 32226 37042
rect 32226 36990 32228 37042
rect 32172 36988 32228 36990
rect 31948 35698 32004 35700
rect 31948 35646 31950 35698
rect 31950 35646 32002 35698
rect 32002 35646 32004 35698
rect 31948 35644 32004 35646
rect 36988 37212 37044 37268
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 40684 42700 40740 42756
rect 42028 45612 42084 45668
rect 41804 45276 41860 45332
rect 42028 45388 42084 45444
rect 41580 45106 41636 45108
rect 41580 45054 41582 45106
rect 41582 45054 41634 45106
rect 41634 45054 41636 45106
rect 41580 45052 41636 45054
rect 41804 44994 41860 44996
rect 41804 44942 41806 44994
rect 41806 44942 41858 44994
rect 41858 44942 41860 44994
rect 41804 44940 41860 44942
rect 42476 48076 42532 48132
rect 42364 46674 42420 46676
rect 42364 46622 42366 46674
rect 42366 46622 42418 46674
rect 42418 46622 42420 46674
rect 42364 46620 42420 46622
rect 42364 45612 42420 45668
rect 42812 49810 42868 49812
rect 42812 49758 42814 49810
rect 42814 49758 42866 49810
rect 42866 49758 42868 49810
rect 42812 49756 42868 49758
rect 44044 49868 44100 49924
rect 43260 49644 43316 49700
rect 43932 49756 43988 49812
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 46620 49980 46676 50036
rect 47628 50034 47684 50036
rect 47628 49982 47630 50034
rect 47630 49982 47682 50034
rect 47682 49982 47684 50034
rect 47628 49980 47684 49982
rect 47740 49922 47796 49924
rect 47740 49870 47742 49922
rect 47742 49870 47794 49922
rect 47794 49870 47796 49922
rect 47740 49868 47796 49870
rect 45948 49756 46004 49812
rect 46956 49810 47012 49812
rect 46956 49758 46958 49810
rect 46958 49758 47010 49810
rect 47010 49758 47012 49810
rect 46956 49756 47012 49758
rect 44044 49698 44100 49700
rect 44044 49646 44046 49698
rect 44046 49646 44098 49698
rect 44098 49646 44100 49698
rect 44044 49644 44100 49646
rect 42700 47068 42756 47124
rect 43036 48076 43092 48132
rect 42700 46620 42756 46676
rect 42588 46450 42644 46452
rect 42588 46398 42590 46450
rect 42590 46398 42642 46450
rect 42642 46398 42644 46450
rect 42588 46396 42644 46398
rect 42140 43538 42196 43540
rect 42140 43486 42142 43538
rect 42142 43486 42194 43538
rect 42194 43486 42196 43538
rect 42140 43484 42196 43486
rect 42476 43484 42532 43540
rect 41580 42866 41636 42868
rect 41580 42814 41582 42866
rect 41582 42814 41634 42866
rect 41634 42814 41636 42866
rect 41580 42812 41636 42814
rect 42364 42866 42420 42868
rect 42364 42814 42366 42866
rect 42366 42814 42418 42866
rect 42418 42814 42420 42866
rect 42364 42812 42420 42814
rect 42252 42754 42308 42756
rect 42252 42702 42254 42754
rect 42254 42702 42306 42754
rect 42306 42702 42308 42754
rect 42252 42700 42308 42702
rect 44716 48860 44772 48916
rect 45500 48914 45556 48916
rect 45500 48862 45502 48914
rect 45502 48862 45554 48914
rect 45554 48862 45556 48914
rect 45500 48860 45556 48862
rect 43708 48076 43764 48132
rect 44492 48130 44548 48132
rect 44492 48078 44494 48130
rect 44494 48078 44546 48130
rect 44546 48078 44548 48130
rect 44492 48076 44548 48078
rect 44492 47292 44548 47348
rect 45612 47346 45668 47348
rect 45612 47294 45614 47346
rect 45614 47294 45666 47346
rect 45666 47294 45668 47346
rect 45612 47292 45668 47294
rect 48972 49756 49028 49812
rect 52444 51266 52500 51268
rect 52444 51214 52446 51266
rect 52446 51214 52498 51266
rect 52498 51214 52500 51266
rect 52444 51212 52500 51214
rect 55132 51212 55188 51268
rect 53340 50428 53396 50484
rect 54236 50482 54292 50484
rect 54236 50430 54238 50482
rect 54238 50430 54290 50482
rect 54290 50430 54292 50482
rect 54236 50428 54292 50430
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 49532 49756 49588 49812
rect 45836 47180 45892 47236
rect 47180 47180 47236 47236
rect 51100 49810 51156 49812
rect 51100 49758 51102 49810
rect 51102 49758 51154 49810
rect 51154 49758 51156 49810
rect 51100 49756 51156 49758
rect 53004 49756 53060 49812
rect 53564 49756 53620 49812
rect 48972 48914 49028 48916
rect 48972 48862 48974 48914
rect 48974 48862 49026 48914
rect 49026 48862 49028 48914
rect 48972 48860 49028 48862
rect 50316 48914 50372 48916
rect 50316 48862 50318 48914
rect 50318 48862 50370 48914
rect 50370 48862 50372 48914
rect 50316 48860 50372 48862
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 48748 48242 48804 48244
rect 48748 48190 48750 48242
rect 48750 48190 48802 48242
rect 48802 48190 48804 48242
rect 48748 48188 48804 48190
rect 49532 48242 49588 48244
rect 49532 48190 49534 48242
rect 49534 48190 49586 48242
rect 49586 48190 49588 48242
rect 49532 48188 49588 48190
rect 50876 48188 50932 48244
rect 50092 47570 50148 47572
rect 50092 47518 50094 47570
rect 50094 47518 50146 47570
rect 50146 47518 50148 47570
rect 50092 47516 50148 47518
rect 47516 47180 47572 47236
rect 48412 46732 48468 46788
rect 43820 45836 43876 45892
rect 47740 46508 47796 46564
rect 47068 46396 47124 46452
rect 46956 45948 47012 46004
rect 43932 45388 43988 45444
rect 46620 44994 46676 44996
rect 46620 44942 46622 44994
rect 46622 44942 46674 44994
rect 46674 44942 46676 44994
rect 46620 44940 46676 44942
rect 47404 44940 47460 44996
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50428 46620 50484 46676
rect 49532 46562 49588 46564
rect 49532 46510 49534 46562
rect 49534 46510 49586 46562
rect 49586 46510 49588 46562
rect 49532 46508 49588 46510
rect 48972 46002 49028 46004
rect 48972 45950 48974 46002
rect 48974 45950 49026 46002
rect 49026 45950 49028 46002
rect 48972 45948 49028 45950
rect 50428 45948 50484 46004
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 48412 44156 48468 44212
rect 48972 44210 49028 44212
rect 48972 44158 48974 44210
rect 48974 44158 49026 44210
rect 49026 44158 49028 44210
rect 48972 44156 49028 44158
rect 48412 43762 48468 43764
rect 48412 43710 48414 43762
rect 48414 43710 48466 43762
rect 48466 43710 48468 43762
rect 48412 43708 48468 43710
rect 43820 42700 43876 42756
rect 44716 42754 44772 42756
rect 44716 42702 44718 42754
rect 44718 42702 44770 42754
rect 44770 42702 44772 42754
rect 44716 42700 44772 42702
rect 44940 42700 44996 42756
rect 42812 42588 42868 42644
rect 44492 42588 44548 42644
rect 42588 42028 42644 42084
rect 45612 42754 45668 42756
rect 45612 42702 45614 42754
rect 45614 42702 45666 42754
rect 45666 42702 45668 42754
rect 45612 42700 45668 42702
rect 49420 43426 49476 43428
rect 49420 43374 49422 43426
rect 49422 43374 49474 43426
rect 49474 43374 49476 43426
rect 49420 43372 49476 43374
rect 46956 42700 47012 42756
rect 54348 48914 54404 48916
rect 54348 48862 54350 48914
rect 54350 48862 54402 48914
rect 54402 48862 54404 48914
rect 54348 48860 54404 48862
rect 52444 47404 52500 47460
rect 53452 47516 53508 47572
rect 54012 47458 54068 47460
rect 54012 47406 54014 47458
rect 54014 47406 54066 47458
rect 54066 47406 54068 47458
rect 54012 47404 54068 47406
rect 52668 47068 52724 47124
rect 51548 46956 51604 47012
rect 51212 46674 51268 46676
rect 51212 46622 51214 46674
rect 51214 46622 51266 46674
rect 51266 46622 51268 46674
rect 51212 46620 51268 46622
rect 54012 46732 54068 46788
rect 51548 46620 51604 46676
rect 55356 49084 55412 49140
rect 56924 48914 56980 48916
rect 56924 48862 56926 48914
rect 56926 48862 56978 48914
rect 56978 48862 56980 48914
rect 56924 48860 56980 48862
rect 54572 46956 54628 47012
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 52444 44268 52500 44324
rect 50876 43372 50932 43428
rect 51100 43708 51156 43764
rect 52332 43596 52388 43652
rect 51212 43372 51268 43428
rect 50876 42700 50932 42756
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 49644 42028 49700 42084
rect 50092 42028 50148 42084
rect 50876 42028 50932 42084
rect 42476 40908 42532 40964
rect 44380 40962 44436 40964
rect 44380 40910 44382 40962
rect 44382 40910 44434 40962
rect 44434 40910 44436 40962
rect 44380 40908 44436 40910
rect 46844 40908 46900 40964
rect 40908 40348 40964 40404
rect 43372 39058 43428 39060
rect 43372 39006 43374 39058
rect 43374 39006 43426 39058
rect 43426 39006 43428 39058
rect 43372 39004 43428 39006
rect 44044 39058 44100 39060
rect 44044 39006 44046 39058
rect 44046 39006 44098 39058
rect 44098 39006 44100 39058
rect 44044 39004 44100 39006
rect 40012 38780 40068 38836
rect 40348 38668 40404 38724
rect 37660 38556 37716 38612
rect 39676 38556 39732 38612
rect 37548 38162 37604 38164
rect 37548 38110 37550 38162
rect 37550 38110 37602 38162
rect 37602 38110 37604 38162
rect 37548 38108 37604 38110
rect 42812 38668 42868 38724
rect 37884 37884 37940 37940
rect 37436 37100 37492 37156
rect 36988 36540 37044 36596
rect 37548 36594 37604 36596
rect 37548 36542 37550 36594
rect 37550 36542 37602 36594
rect 37602 36542 37604 36594
rect 37548 36540 37604 36542
rect 33068 35532 33124 35588
rect 36092 35586 36148 35588
rect 36092 35534 36094 35586
rect 36094 35534 36146 35586
rect 36146 35534 36148 35586
rect 36092 35532 36148 35534
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35308 34018 35364 34020
rect 35308 33966 35310 34018
rect 35310 33966 35362 34018
rect 35362 33966 35364 34018
rect 35308 33964 35364 33966
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 27020 32396 27076 32452
rect 24108 29372 24164 29428
rect 24892 28812 24948 28868
rect 25900 28866 25956 28868
rect 25900 28814 25902 28866
rect 25902 28814 25954 28866
rect 25954 28814 25956 28866
rect 25900 28812 25956 28814
rect 21196 28364 21252 28420
rect 16380 27746 16436 27748
rect 16380 27694 16382 27746
rect 16382 27694 16434 27746
rect 16434 27694 16436 27746
rect 16380 27692 16436 27694
rect 15820 27244 15876 27300
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 15820 25506 15876 25508
rect 15820 25454 15822 25506
rect 15822 25454 15874 25506
rect 15874 25454 15876 25506
rect 15820 25452 15876 25454
rect 21756 28082 21812 28084
rect 21756 28030 21758 28082
rect 21758 28030 21810 28082
rect 21810 28030 21812 28082
rect 21756 28028 21812 28030
rect 21532 27916 21588 27972
rect 18620 25618 18676 25620
rect 18620 25566 18622 25618
rect 18622 25566 18674 25618
rect 18674 25566 18676 25618
rect 18620 25564 18676 25566
rect 20300 25618 20356 25620
rect 20300 25566 20302 25618
rect 20302 25566 20354 25618
rect 20354 25566 20356 25618
rect 20300 25564 20356 25566
rect 17836 25452 17892 25508
rect 18284 25452 18340 25508
rect 16492 24892 16548 24948
rect 17724 24946 17780 24948
rect 17724 24894 17726 24946
rect 17726 24894 17778 24946
rect 17778 24894 17780 24946
rect 17724 24892 17780 24894
rect 20188 25506 20244 25508
rect 20188 25454 20190 25506
rect 20190 25454 20242 25506
rect 20242 25454 20244 25506
rect 20188 25452 20244 25454
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 17052 24050 17108 24052
rect 17052 23998 17054 24050
rect 17054 23998 17106 24050
rect 17106 23998 17108 24050
rect 17052 23996 17108 23998
rect 16604 23548 16660 23604
rect 17948 23660 18004 23716
rect 16604 23378 16660 23380
rect 16604 23326 16606 23378
rect 16606 23326 16658 23378
rect 16658 23326 16660 23378
rect 16604 23324 16660 23326
rect 15260 22482 15316 22484
rect 15260 22430 15262 22482
rect 15262 22430 15314 22482
rect 15314 22430 15316 22482
rect 15260 22428 15316 22430
rect 13132 21532 13188 21588
rect 13468 20524 13524 20580
rect 12572 19346 12628 19348
rect 12572 19294 12574 19346
rect 12574 19294 12626 19346
rect 12626 19294 12628 19346
rect 12572 19292 12628 19294
rect 11788 17724 11844 17780
rect 9660 16828 9716 16884
rect 8764 16716 8820 16772
rect 10780 16882 10836 16884
rect 10780 16830 10782 16882
rect 10782 16830 10834 16882
rect 10834 16830 10836 16882
rect 10780 16828 10836 16830
rect 11452 16882 11508 16884
rect 11452 16830 11454 16882
rect 11454 16830 11506 16882
rect 11506 16830 11508 16882
rect 11452 16828 11508 16830
rect 11564 16210 11620 16212
rect 11564 16158 11566 16210
rect 11566 16158 11618 16210
rect 11618 16158 11620 16210
rect 11564 16156 11620 16158
rect 8764 15036 8820 15092
rect 8652 13692 8708 13748
rect 8988 13804 9044 13860
rect 8988 12962 9044 12964
rect 8988 12910 8990 12962
rect 8990 12910 9042 12962
rect 9042 12910 9044 12962
rect 8988 12908 9044 12910
rect 9100 12850 9156 12852
rect 9100 12798 9102 12850
rect 9102 12798 9154 12850
rect 9154 12798 9156 12850
rect 9100 12796 9156 12798
rect 11340 15036 11396 15092
rect 9996 13746 10052 13748
rect 9996 13694 9998 13746
rect 9998 13694 10050 13746
rect 10050 13694 10052 13746
rect 9996 13692 10052 13694
rect 8316 12124 8372 12180
rect 8988 12178 9044 12180
rect 8988 12126 8990 12178
rect 8990 12126 9042 12178
rect 9042 12126 9044 12178
rect 8988 12124 9044 12126
rect 8204 11340 8260 11396
rect 7308 10556 7364 10612
rect 3948 10498 4004 10500
rect 3948 10446 3950 10498
rect 3950 10446 4002 10498
rect 4002 10446 4004 10498
rect 3948 10444 4004 10446
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 7196 9884 7252 9940
rect 6972 9826 7028 9828
rect 6972 9774 6974 9826
rect 6974 9774 7026 9826
rect 7026 9774 7028 9826
rect 6972 9772 7028 9774
rect 4732 9660 4788 9716
rect 3388 9100 3444 9156
rect 4060 9042 4116 9044
rect 4060 8990 4062 9042
rect 4062 8990 4114 9042
rect 4114 8990 4116 9042
rect 4060 8988 4116 8990
rect 6748 9714 6804 9716
rect 6748 9662 6750 9714
rect 6750 9662 6802 9714
rect 6802 9662 6804 9714
rect 6748 9660 6804 9662
rect 6860 9436 6916 9492
rect 5964 9154 6020 9156
rect 5964 9102 5966 9154
rect 5966 9102 6018 9154
rect 6018 9102 6020 9154
rect 5964 9100 6020 9102
rect 6860 9100 6916 9156
rect 7196 9660 7252 9716
rect 4732 8988 4788 9044
rect 4956 8988 5012 9044
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 6188 9042 6244 9044
rect 6188 8990 6190 9042
rect 6190 8990 6242 9042
rect 6242 8990 6244 9042
rect 6188 8988 6244 8990
rect 8204 10556 8260 10612
rect 8092 9938 8148 9940
rect 8092 9886 8094 9938
rect 8094 9886 8146 9938
rect 8146 9886 8148 9938
rect 8092 9884 8148 9886
rect 7420 9602 7476 9604
rect 7420 9550 7422 9602
rect 7422 9550 7474 9602
rect 7474 9550 7476 9602
rect 7420 9548 7476 9550
rect 7868 9436 7924 9492
rect 9772 12402 9828 12404
rect 9772 12350 9774 12402
rect 9774 12350 9826 12402
rect 9826 12350 9828 12402
rect 9772 12348 9828 12350
rect 9548 11900 9604 11956
rect 10108 11954 10164 11956
rect 10108 11902 10110 11954
rect 10110 11902 10162 11954
rect 10162 11902 10164 11954
rect 10108 11900 10164 11902
rect 10444 13746 10500 13748
rect 10444 13694 10446 13746
rect 10446 13694 10498 13746
rect 10498 13694 10500 13746
rect 10444 13692 10500 13694
rect 13132 18172 13188 18228
rect 13916 19292 13972 19348
rect 12796 16716 12852 16772
rect 13580 17778 13636 17780
rect 13580 17726 13582 17778
rect 13582 17726 13634 17778
rect 13634 17726 13636 17778
rect 13580 17724 13636 17726
rect 14140 18450 14196 18452
rect 14140 18398 14142 18450
rect 14142 18398 14194 18450
rect 14194 18398 14196 18450
rect 14140 18396 14196 18398
rect 14812 18338 14868 18340
rect 14812 18286 14814 18338
rect 14814 18286 14866 18338
rect 14866 18286 14868 18338
rect 14812 18284 14868 18286
rect 16044 22428 16100 22484
rect 17388 22482 17444 22484
rect 17388 22430 17390 22482
rect 17390 22430 17442 22482
rect 17442 22430 17444 22482
rect 17388 22428 17444 22430
rect 18284 23660 18340 23716
rect 20748 24556 20804 24612
rect 20860 25452 20916 25508
rect 18844 23660 18900 23716
rect 18508 23548 18564 23604
rect 18060 22428 18116 22484
rect 16828 19906 16884 19908
rect 16828 19854 16830 19906
rect 16830 19854 16882 19906
rect 16882 19854 16884 19906
rect 16828 19852 16884 19854
rect 15596 19292 15652 19348
rect 16940 19740 16996 19796
rect 15484 18284 15540 18340
rect 16604 18396 16660 18452
rect 13804 16210 13860 16212
rect 13804 16158 13806 16210
rect 13806 16158 13858 16210
rect 13858 16158 13860 16210
rect 13804 16156 13860 16158
rect 13132 15202 13188 15204
rect 13132 15150 13134 15202
rect 13134 15150 13186 15202
rect 13186 15150 13188 15202
rect 13132 15148 13188 15150
rect 20188 23660 20244 23716
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18732 20188 18788 20244
rect 18284 19906 18340 19908
rect 18284 19854 18286 19906
rect 18286 19854 18338 19906
rect 18338 19854 18340 19906
rect 18284 19852 18340 19854
rect 17052 18284 17108 18340
rect 17276 18284 17332 18340
rect 17836 19794 17892 19796
rect 17836 19742 17838 19794
rect 17838 19742 17890 19794
rect 17890 19742 17892 19794
rect 17836 19740 17892 19742
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 25004 27858 25060 27860
rect 25004 27806 25006 27858
rect 25006 27806 25058 27858
rect 25058 27806 25060 27858
rect 25004 27804 25060 27806
rect 25788 28418 25844 28420
rect 25788 28366 25790 28418
rect 25790 28366 25842 28418
rect 25842 28366 25844 28418
rect 25788 28364 25844 28366
rect 25676 27858 25732 27860
rect 25676 27806 25678 27858
rect 25678 27806 25730 27858
rect 25730 27806 25732 27858
rect 25676 27804 25732 27806
rect 23996 26460 24052 26516
rect 21644 25452 21700 25508
rect 22316 25506 22372 25508
rect 22316 25454 22318 25506
rect 22318 25454 22370 25506
rect 22370 25454 22372 25506
rect 22316 25452 22372 25454
rect 24892 26514 24948 26516
rect 24892 26462 24894 26514
rect 24894 26462 24946 26514
rect 24946 26462 24948 26514
rect 24892 26460 24948 26462
rect 25564 26460 25620 26516
rect 24444 26178 24500 26180
rect 24444 26126 24446 26178
rect 24446 26126 24498 26178
rect 24498 26126 24500 26178
rect 24444 26124 24500 26126
rect 25116 25618 25172 25620
rect 25116 25566 25118 25618
rect 25118 25566 25170 25618
rect 25170 25566 25172 25618
rect 25116 25564 25172 25566
rect 27244 29932 27300 29988
rect 26572 29426 26628 29428
rect 26572 29374 26574 29426
rect 26574 29374 26626 29426
rect 26626 29374 26628 29426
rect 26572 29372 26628 29374
rect 32732 32620 32788 32676
rect 31948 31500 32004 31556
rect 29708 30994 29764 30996
rect 29708 30942 29710 30994
rect 29710 30942 29762 30994
rect 29762 30942 29764 30994
rect 29708 30940 29764 30942
rect 29932 30940 29988 30996
rect 28140 29986 28196 29988
rect 28140 29934 28142 29986
rect 28142 29934 28194 29986
rect 28194 29934 28196 29986
rect 28140 29932 28196 29934
rect 27356 29372 27412 29428
rect 28140 29372 28196 29428
rect 26348 28028 26404 28084
rect 27692 28028 27748 28084
rect 26236 27916 26292 27972
rect 26124 26124 26180 26180
rect 26348 27804 26404 27860
rect 25788 25564 25844 25620
rect 23996 25452 24052 25508
rect 21756 24610 21812 24612
rect 21756 24558 21758 24610
rect 21758 24558 21810 24610
rect 21810 24558 21812 24610
rect 21756 24556 21812 24558
rect 20972 23660 21028 23716
rect 24668 24050 24724 24052
rect 24668 23998 24670 24050
rect 24670 23998 24722 24050
rect 24722 23998 24724 24050
rect 24668 23996 24724 23998
rect 25676 23996 25732 24052
rect 22204 23660 22260 23716
rect 33628 32674 33684 32676
rect 33628 32622 33630 32674
rect 33630 32622 33682 32674
rect 33682 32622 33684 32674
rect 33628 32620 33684 32622
rect 36540 34188 36596 34244
rect 37436 34242 37492 34244
rect 37436 34190 37438 34242
rect 37438 34190 37490 34242
rect 37490 34190 37492 34242
rect 37436 34188 37492 34190
rect 36428 33964 36484 34020
rect 36316 33068 36372 33124
rect 36540 33292 36596 33348
rect 38332 37490 38388 37492
rect 38332 37438 38334 37490
rect 38334 37438 38386 37490
rect 38386 37438 38388 37490
rect 38332 37436 38388 37438
rect 40796 36428 40852 36484
rect 39452 35196 39508 35252
rect 38220 34130 38276 34132
rect 38220 34078 38222 34130
rect 38222 34078 38274 34130
rect 38274 34078 38276 34130
rect 38220 34076 38276 34078
rect 39452 34076 39508 34132
rect 40572 35196 40628 35252
rect 37660 33292 37716 33348
rect 42924 37436 42980 37492
rect 43484 38834 43540 38836
rect 43484 38782 43486 38834
rect 43486 38782 43538 38834
rect 43538 38782 43540 38834
rect 43484 38780 43540 38782
rect 46620 39676 46676 39732
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 47628 39730 47684 39732
rect 47628 39678 47630 39730
rect 47630 39678 47682 39730
rect 47682 39678 47684 39730
rect 47628 39676 47684 39678
rect 46844 39564 46900 39620
rect 44380 38722 44436 38724
rect 44380 38670 44382 38722
rect 44382 38670 44434 38722
rect 44434 38670 44436 38722
rect 44380 38668 44436 38670
rect 43484 36540 43540 36596
rect 43148 36482 43204 36484
rect 43148 36430 43150 36482
rect 43150 36430 43202 36482
rect 43202 36430 43204 36482
rect 43148 36428 43204 36430
rect 41468 35196 41524 35252
rect 41804 35308 41860 35364
rect 40572 33628 40628 33684
rect 41356 34076 41412 34132
rect 36764 33122 36820 33124
rect 36764 33070 36766 33122
rect 36766 33070 36818 33122
rect 36818 33070 36820 33122
rect 36764 33068 36820 33070
rect 37660 33068 37716 33124
rect 34748 32284 34804 32340
rect 35980 32338 36036 32340
rect 35980 32286 35982 32338
rect 35982 32286 36034 32338
rect 36034 32286 36036 32338
rect 35980 32284 36036 32286
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 32508 31500 32564 31556
rect 33740 31500 33796 31556
rect 35196 31554 35252 31556
rect 35196 31502 35198 31554
rect 35198 31502 35250 31554
rect 35250 31502 35252 31554
rect 35196 31500 35252 31502
rect 31948 30940 32004 30996
rect 32284 30322 32340 30324
rect 32284 30270 32286 30322
rect 32286 30270 32338 30322
rect 32338 30270 32340 30322
rect 32284 30268 32340 30270
rect 28252 28642 28308 28644
rect 28252 28590 28254 28642
rect 28254 28590 28306 28642
rect 28306 28590 28308 28642
rect 28252 28588 28308 28590
rect 28140 26460 28196 26516
rect 26796 24050 26852 24052
rect 26796 23998 26798 24050
rect 26798 23998 26850 24050
rect 26850 23998 26852 24050
rect 26796 23996 26852 23998
rect 23436 23266 23492 23268
rect 23436 23214 23438 23266
rect 23438 23214 23490 23266
rect 23490 23214 23492 23266
rect 23436 23212 23492 23214
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19516 20242 19572 20244
rect 19516 20190 19518 20242
rect 19518 20190 19570 20242
rect 19570 20190 19572 20242
rect 19516 20188 19572 20190
rect 23212 21644 23268 21700
rect 20860 20914 20916 20916
rect 20860 20862 20862 20914
rect 20862 20862 20914 20914
rect 20914 20862 20916 20914
rect 20860 20860 20916 20862
rect 19180 19068 19236 19124
rect 19516 19068 19572 19124
rect 19404 18508 19460 18564
rect 17948 18450 18004 18452
rect 17948 18398 17950 18450
rect 17950 18398 18002 18450
rect 18002 18398 18004 18450
rect 17948 18396 18004 18398
rect 17724 18172 17780 18228
rect 19292 16828 19348 16884
rect 20076 19122 20132 19124
rect 20076 19070 20078 19122
rect 20078 19070 20130 19122
rect 20130 19070 20132 19122
rect 20076 19068 20132 19070
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 22540 19852 22596 19908
rect 21532 19346 21588 19348
rect 21532 19294 21534 19346
rect 21534 19294 21586 19346
rect 21586 19294 21588 19346
rect 21532 19292 21588 19294
rect 21196 18508 21252 18564
rect 26348 23212 26404 23268
rect 26684 23660 26740 23716
rect 22988 19068 23044 19124
rect 27356 23714 27412 23716
rect 27356 23662 27358 23714
rect 27358 23662 27410 23714
rect 27410 23662 27412 23714
rect 27356 23660 27412 23662
rect 26908 23154 26964 23156
rect 26908 23102 26910 23154
rect 26910 23102 26962 23154
rect 26962 23102 26964 23154
rect 26908 23100 26964 23102
rect 26012 22370 26068 22372
rect 26012 22318 26014 22370
rect 26014 22318 26066 22370
rect 26066 22318 26068 22370
rect 26012 22316 26068 22318
rect 25676 21698 25732 21700
rect 25676 21646 25678 21698
rect 25678 21646 25730 21698
rect 25730 21646 25732 21698
rect 25676 21644 25732 21646
rect 24332 20860 24388 20916
rect 24556 20860 24612 20916
rect 25340 20914 25396 20916
rect 25340 20862 25342 20914
rect 25342 20862 25394 20914
rect 25394 20862 25396 20914
rect 25340 20860 25396 20862
rect 26684 20188 26740 20244
rect 24556 19906 24612 19908
rect 24556 19854 24558 19906
rect 24558 19854 24610 19906
rect 24610 19854 24612 19906
rect 24556 19852 24612 19854
rect 25452 19852 25508 19908
rect 22540 18508 22596 18564
rect 22764 18508 22820 18564
rect 19516 17836 19572 17892
rect 14364 15148 14420 15204
rect 18844 15314 18900 15316
rect 18844 15262 18846 15314
rect 18846 15262 18898 15314
rect 18898 15262 18900 15314
rect 18844 15260 18900 15262
rect 19628 18396 19684 18452
rect 21308 18450 21364 18452
rect 21308 18398 21310 18450
rect 21310 18398 21362 18450
rect 21362 18398 21364 18450
rect 21308 18396 21364 18398
rect 20748 18338 20804 18340
rect 20748 18286 20750 18338
rect 20750 18286 20802 18338
rect 20802 18286 20804 18338
rect 20748 18284 20804 18286
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 21980 18338 22036 18340
rect 21980 18286 21982 18338
rect 21982 18286 22034 18338
rect 22034 18286 22036 18338
rect 21980 18284 22036 18286
rect 21756 16828 21812 16884
rect 22540 18226 22596 18228
rect 22540 18174 22542 18226
rect 22542 18174 22594 18226
rect 22594 18174 22596 18226
rect 22540 18172 22596 18174
rect 23324 18172 23380 18228
rect 25788 17106 25844 17108
rect 25788 17054 25790 17106
rect 25790 17054 25842 17106
rect 25842 17054 25844 17106
rect 25788 17052 25844 17054
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19516 15314 19572 15316
rect 19516 15262 19518 15314
rect 19518 15262 19570 15314
rect 19570 15262 19572 15314
rect 19516 15260 19572 15262
rect 22540 15820 22596 15876
rect 20188 15036 20244 15092
rect 16268 14306 16324 14308
rect 16268 14254 16270 14306
rect 16270 14254 16322 14306
rect 16322 14254 16324 14306
rect 16268 14252 16324 14254
rect 16828 14252 16884 14308
rect 17276 14252 17332 14308
rect 12572 13692 12628 13748
rect 10668 12962 10724 12964
rect 10668 12910 10670 12962
rect 10670 12910 10722 12962
rect 10722 12910 10724 12962
rect 10668 12908 10724 12910
rect 10332 12796 10388 12852
rect 8540 9826 8596 9828
rect 8540 9774 8542 9826
rect 8542 9774 8594 9826
rect 8594 9774 8596 9826
rect 8540 9772 8596 9774
rect 8316 9714 8372 9716
rect 8316 9662 8318 9714
rect 8318 9662 8370 9714
rect 8370 9662 8372 9714
rect 8316 9660 8372 9662
rect 7644 9154 7700 9156
rect 7644 9102 7646 9154
rect 7646 9102 7698 9154
rect 7698 9102 7700 9154
rect 7644 9100 7700 9102
rect 7420 9042 7476 9044
rect 7420 8990 7422 9042
rect 7422 8990 7474 9042
rect 7474 8990 7476 9042
rect 7420 8988 7476 8990
rect 7980 9042 8036 9044
rect 7980 8990 7982 9042
rect 7982 8990 8034 9042
rect 8034 8990 8036 9042
rect 7980 8988 8036 8990
rect 8652 9548 8708 9604
rect 8876 9154 8932 9156
rect 8876 9102 8878 9154
rect 8878 9102 8930 9154
rect 8930 9102 8932 9154
rect 8876 9100 8932 9102
rect 8540 8988 8596 9044
rect 8988 8818 9044 8820
rect 8988 8766 8990 8818
rect 8990 8766 9042 8818
rect 9042 8766 9044 8818
rect 8988 8764 9044 8766
rect 6524 8370 6580 8372
rect 6524 8318 6526 8370
rect 6526 8318 6578 8370
rect 6578 8318 6580 8370
rect 6524 8316 6580 8318
rect 3948 7586 4004 7588
rect 3948 7534 3950 7586
rect 3950 7534 4002 7586
rect 4002 7534 4004 7586
rect 3948 7532 4004 7534
rect 4844 7532 4900 7588
rect 2604 7474 2660 7476
rect 2604 7422 2606 7474
rect 2606 7422 2658 7474
rect 2658 7422 2660 7474
rect 2604 7420 2660 7422
rect 3724 7420 3780 7476
rect 2268 6690 2324 6692
rect 2268 6638 2270 6690
rect 2270 6638 2322 6690
rect 2322 6638 2324 6690
rect 2268 6636 2324 6638
rect 2716 6690 2772 6692
rect 2716 6638 2718 6690
rect 2718 6638 2770 6690
rect 2770 6638 2772 6690
rect 2716 6636 2772 6638
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4172 6690 4228 6692
rect 4172 6638 4174 6690
rect 4174 6638 4226 6690
rect 4226 6638 4228 6690
rect 4172 6636 4228 6638
rect 3724 6578 3780 6580
rect 3724 6526 3726 6578
rect 3726 6526 3778 6578
rect 3778 6526 3780 6578
rect 3724 6524 3780 6526
rect 2828 5964 2884 6020
rect 3948 6018 4004 6020
rect 3948 5966 3950 6018
rect 3950 5966 4002 6018
rect 4002 5966 4004 6018
rect 3948 5964 4004 5966
rect 9772 10444 9828 10500
rect 10220 11340 10276 11396
rect 10668 11170 10724 11172
rect 10668 11118 10670 11170
rect 10670 11118 10722 11170
rect 10722 11118 10724 11170
rect 10668 11116 10724 11118
rect 11004 12738 11060 12740
rect 11004 12686 11006 12738
rect 11006 12686 11058 12738
rect 11058 12686 11060 12738
rect 11004 12684 11060 12686
rect 11004 12178 11060 12180
rect 11004 12126 11006 12178
rect 11006 12126 11058 12178
rect 11058 12126 11060 12178
rect 11004 12124 11060 12126
rect 12572 12962 12628 12964
rect 12572 12910 12574 12962
rect 12574 12910 12626 12962
rect 12626 12910 12628 12962
rect 12572 12908 12628 12910
rect 11340 12850 11396 12852
rect 11340 12798 11342 12850
rect 11342 12798 11394 12850
rect 11394 12798 11396 12850
rect 11340 12796 11396 12798
rect 11900 12850 11956 12852
rect 11900 12798 11902 12850
rect 11902 12798 11954 12850
rect 11954 12798 11956 12850
rect 11900 12796 11956 12798
rect 11676 12684 11732 12740
rect 11116 11900 11172 11956
rect 12124 11788 12180 11844
rect 11004 11116 11060 11172
rect 9884 10108 9940 10164
rect 5740 7532 5796 7588
rect 8540 7532 8596 7588
rect 9324 9602 9380 9604
rect 9324 9550 9326 9602
rect 9326 9550 9378 9602
rect 9378 9550 9380 9602
rect 9324 9548 9380 9550
rect 9996 10444 10052 10500
rect 10220 9602 10276 9604
rect 10220 9550 10222 9602
rect 10222 9550 10274 9602
rect 10274 9550 10276 9602
rect 10220 9548 10276 9550
rect 11900 11170 11956 11172
rect 11900 11118 11902 11170
rect 11902 11118 11954 11170
rect 11954 11118 11956 11170
rect 11900 11116 11956 11118
rect 11004 10610 11060 10612
rect 11004 10558 11006 10610
rect 11006 10558 11058 10610
rect 11058 10558 11060 10610
rect 11004 10556 11060 10558
rect 13804 12908 13860 12964
rect 13356 12684 13412 12740
rect 13356 12124 13412 12180
rect 13020 11788 13076 11844
rect 12236 11116 12292 11172
rect 11228 10108 11284 10164
rect 10780 9548 10836 9604
rect 10220 8818 10276 8820
rect 10220 8766 10222 8818
rect 10222 8766 10274 8818
rect 10274 8766 10276 8818
rect 10220 8764 10276 8766
rect 11004 9100 11060 9156
rect 10108 8316 10164 8372
rect 10108 8146 10164 8148
rect 10108 8094 10110 8146
rect 10110 8094 10162 8146
rect 10162 8094 10164 8146
rect 10108 8092 10164 8094
rect 11340 9714 11396 9716
rect 11340 9662 11342 9714
rect 11342 9662 11394 9714
rect 11394 9662 11396 9714
rect 11340 9660 11396 9662
rect 11900 9714 11956 9716
rect 11900 9662 11902 9714
rect 11902 9662 11954 9714
rect 11954 9662 11956 9714
rect 11900 9660 11956 9662
rect 12684 11170 12740 11172
rect 12684 11118 12686 11170
rect 12686 11118 12738 11170
rect 12738 11118 12740 11170
rect 12684 11116 12740 11118
rect 12572 9826 12628 9828
rect 12572 9774 12574 9826
rect 12574 9774 12626 9826
rect 12626 9774 12628 9826
rect 12572 9772 12628 9774
rect 12796 9042 12852 9044
rect 12796 8990 12798 9042
rect 12798 8990 12850 9042
rect 12850 8990 12852 9042
rect 12796 8988 12852 8990
rect 16940 13132 16996 13188
rect 14812 12796 14868 12852
rect 15596 12850 15652 12852
rect 15596 12798 15598 12850
rect 15598 12798 15650 12850
rect 15650 12798 15652 12850
rect 15596 12796 15652 12798
rect 14028 12738 14084 12740
rect 14028 12686 14030 12738
rect 14030 12686 14082 12738
rect 14082 12686 14084 12738
rect 14028 12684 14084 12686
rect 13804 12124 13860 12180
rect 14252 11954 14308 11956
rect 14252 11902 14254 11954
rect 14254 11902 14306 11954
rect 14306 11902 14308 11954
rect 14252 11900 14308 11902
rect 14028 11170 14084 11172
rect 14028 11118 14030 11170
rect 14030 11118 14082 11170
rect 14082 11118 14084 11170
rect 14028 11116 14084 11118
rect 14476 12178 14532 12180
rect 14476 12126 14478 12178
rect 14478 12126 14530 12178
rect 14530 12126 14532 12178
rect 14476 12124 14532 12126
rect 14364 11116 14420 11172
rect 15596 11788 15652 11844
rect 16156 11452 16212 11508
rect 19292 13186 19348 13188
rect 19292 13134 19294 13186
rect 19294 13134 19346 13186
rect 19346 13134 19348 13186
rect 19292 13132 19348 13134
rect 20412 15260 20468 15316
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 15596 9772 15652 9828
rect 13468 9154 13524 9156
rect 13468 9102 13470 9154
rect 13470 9102 13522 9154
rect 13522 9102 13524 9154
rect 13468 9100 13524 9102
rect 13356 8988 13412 9044
rect 15484 8988 15540 9044
rect 11004 8092 11060 8148
rect 10780 7362 10836 7364
rect 10780 7310 10782 7362
rect 10782 7310 10834 7362
rect 10834 7310 10836 7362
rect 10780 7308 10836 7310
rect 11340 6802 11396 6804
rect 11340 6750 11342 6802
rect 11342 6750 11394 6802
rect 11394 6750 11396 6802
rect 11340 6748 11396 6750
rect 11452 7308 11508 7364
rect 9100 6524 9156 6580
rect 12124 7532 12180 7588
rect 14700 7586 14756 7588
rect 14700 7534 14702 7586
rect 14702 7534 14754 7586
rect 14754 7534 14756 7586
rect 14700 7532 14756 7534
rect 15708 8988 15764 9044
rect 16044 9042 16100 9044
rect 16044 8990 16046 9042
rect 16046 8990 16098 9042
rect 16098 8990 16100 9042
rect 16044 8988 16100 8990
rect 16828 9884 16884 9940
rect 19964 13074 20020 13076
rect 19964 13022 19966 13074
rect 19966 13022 20018 13074
rect 20018 13022 20020 13074
rect 19964 13020 20020 13022
rect 16828 8988 16884 9044
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 20636 15036 20692 15092
rect 21420 15036 21476 15092
rect 21756 15036 21812 15092
rect 23772 15874 23828 15876
rect 23772 15822 23774 15874
rect 23774 15822 23826 15874
rect 23826 15822 23828 15874
rect 23772 15820 23828 15822
rect 21756 13916 21812 13972
rect 23884 13970 23940 13972
rect 23884 13918 23886 13970
rect 23886 13918 23938 13970
rect 23938 13918 23940 13970
rect 23884 13916 23940 13918
rect 23324 13074 23380 13076
rect 23324 13022 23326 13074
rect 23326 13022 23378 13074
rect 23378 13022 23380 13074
rect 23324 13020 23380 13022
rect 24668 14642 24724 14644
rect 24668 14590 24670 14642
rect 24670 14590 24722 14642
rect 24722 14590 24724 14642
rect 24668 14588 24724 14590
rect 25564 13468 25620 13524
rect 20412 11506 20468 11508
rect 20412 11454 20414 11506
rect 20414 11454 20466 11506
rect 20466 11454 20468 11506
rect 20412 11452 20468 11454
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19068 9938 19124 9940
rect 19068 9886 19070 9938
rect 19070 9886 19122 9938
rect 19122 9886 19124 9938
rect 19068 9884 19124 9886
rect 19068 9266 19124 9268
rect 19068 9214 19070 9266
rect 19070 9214 19122 9266
rect 19122 9214 19124 9266
rect 19068 9212 19124 9214
rect 12012 7308 12068 7364
rect 12236 6802 12292 6804
rect 12236 6750 12238 6802
rect 12238 6750 12290 6802
rect 12290 6750 12292 6802
rect 12236 6748 12292 6750
rect 11900 6636 11956 6692
rect 19740 10220 19796 10276
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 21980 10556 22036 10612
rect 20412 9212 20468 9268
rect 21868 10220 21924 10276
rect 22204 9826 22260 9828
rect 22204 9774 22206 9826
rect 22206 9774 22258 9826
rect 22258 9774 22260 9826
rect 22204 9772 22260 9774
rect 22092 8482 22148 8484
rect 22092 8430 22094 8482
rect 22094 8430 22146 8482
rect 22146 8430 22148 8482
rect 22092 8428 22148 8430
rect 20860 8258 20916 8260
rect 20860 8206 20862 8258
rect 20862 8206 20914 8258
rect 20914 8206 20916 8258
rect 20860 8204 20916 8206
rect 21868 8258 21924 8260
rect 21868 8206 21870 8258
rect 21870 8206 21922 8258
rect 21922 8206 21924 8258
rect 21868 8204 21924 8206
rect 22652 10610 22708 10612
rect 22652 10558 22654 10610
rect 22654 10558 22706 10610
rect 22706 10558 22708 10610
rect 22652 10556 22708 10558
rect 22988 10498 23044 10500
rect 22988 10446 22990 10498
rect 22990 10446 23042 10498
rect 23042 10446 23044 10498
rect 22988 10444 23044 10446
rect 22428 9772 22484 9828
rect 22876 8482 22932 8484
rect 22876 8430 22878 8482
rect 22878 8430 22930 8482
rect 22930 8430 22932 8482
rect 22876 8428 22932 8430
rect 15820 6636 15876 6692
rect 19180 6636 19236 6692
rect 19628 7980 19684 8036
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20748 8034 20804 8036
rect 20748 7982 20750 8034
rect 20750 7982 20802 8034
rect 20802 7982 20804 8034
rect 20748 7980 20804 7982
rect 20636 7420 20692 7476
rect 22092 7420 22148 7476
rect 19964 7362 20020 7364
rect 19964 7310 19966 7362
rect 19966 7310 20018 7362
rect 20018 7310 20020 7362
rect 19964 7308 20020 7310
rect 22652 7362 22708 7364
rect 22652 7310 22654 7362
rect 22654 7310 22706 7362
rect 22706 7310 22708 7362
rect 22652 7308 22708 7310
rect 24108 12178 24164 12180
rect 24108 12126 24110 12178
rect 24110 12126 24162 12178
rect 24162 12126 24164 12178
rect 24108 12124 24164 12126
rect 23100 7420 23156 7476
rect 22764 7196 22820 7252
rect 22092 6636 22148 6692
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 25004 11618 25060 11620
rect 25004 11566 25006 11618
rect 25006 11566 25058 11618
rect 25058 11566 25060 11618
rect 25004 11564 25060 11566
rect 25452 11564 25508 11620
rect 24668 10444 24724 10500
rect 22092 6076 22148 6132
rect 22428 6130 22484 6132
rect 22428 6078 22430 6130
rect 22430 6078 22482 6130
rect 22482 6078 22484 6130
rect 22428 6076 22484 6078
rect 23212 6076 23268 6132
rect 24668 9826 24724 9828
rect 24668 9774 24670 9826
rect 24670 9774 24722 9826
rect 24722 9774 24724 9826
rect 24668 9772 24724 9774
rect 24892 9826 24948 9828
rect 24892 9774 24894 9826
rect 24894 9774 24946 9826
rect 24946 9774 24948 9826
rect 24892 9772 24948 9774
rect 24668 9212 24724 9268
rect 28588 26460 28644 26516
rect 30268 28642 30324 28644
rect 30268 28590 30270 28642
rect 30270 28590 30322 28642
rect 30322 28590 30324 28642
rect 30268 28588 30324 28590
rect 29372 27804 29428 27860
rect 32732 30322 32788 30324
rect 32732 30270 32734 30322
rect 32734 30270 32786 30322
rect 32786 30270 32788 30322
rect 32732 30268 32788 30270
rect 33292 30322 33348 30324
rect 33292 30270 33294 30322
rect 33294 30270 33346 30322
rect 33346 30270 33348 30322
rect 33292 30268 33348 30270
rect 36764 31052 36820 31108
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 37884 31106 37940 31108
rect 37884 31054 37886 31106
rect 37886 31054 37938 31106
rect 37938 31054 37940 31106
rect 37884 31052 37940 31054
rect 37660 30156 37716 30212
rect 38556 30210 38612 30212
rect 38556 30158 38558 30210
rect 38558 30158 38610 30210
rect 38610 30158 38612 30210
rect 38556 30156 38612 30158
rect 36988 30044 37044 30100
rect 33740 29426 33796 29428
rect 33740 29374 33742 29426
rect 33742 29374 33794 29426
rect 33794 29374 33796 29426
rect 33740 29372 33796 29374
rect 36988 29426 37044 29428
rect 36988 29374 36990 29426
rect 36990 29374 37042 29426
rect 37042 29374 37044 29426
rect 36988 29372 37044 29374
rect 39676 30268 39732 30324
rect 40236 30268 40292 30324
rect 40348 30098 40404 30100
rect 40348 30046 40350 30098
rect 40350 30046 40402 30098
rect 40402 30046 40404 30098
rect 40348 30044 40404 30046
rect 40796 30044 40852 30100
rect 40796 29372 40852 29428
rect 31500 27858 31556 27860
rect 31500 27806 31502 27858
rect 31502 27806 31554 27858
rect 31554 27806 31556 27858
rect 31500 27804 31556 27806
rect 30492 26460 30548 26516
rect 31388 27580 31444 27636
rect 31948 27634 32004 27636
rect 31948 27582 31950 27634
rect 31950 27582 32002 27634
rect 32002 27582 32004 27634
rect 31948 27580 32004 27582
rect 31836 26514 31892 26516
rect 31836 26462 31838 26514
rect 31838 26462 31890 26514
rect 31890 26462 31892 26514
rect 31836 26460 31892 26462
rect 33404 28700 33460 28756
rect 32284 26908 32340 26964
rect 31388 25506 31444 25508
rect 31388 25454 31390 25506
rect 31390 25454 31442 25506
rect 31442 25454 31444 25506
rect 31388 25452 31444 25454
rect 29708 24050 29764 24052
rect 29708 23998 29710 24050
rect 29710 23998 29762 24050
rect 29762 23998 29764 24050
rect 29708 23996 29764 23998
rect 27692 22988 27748 23044
rect 27692 22316 27748 22372
rect 28924 23042 28980 23044
rect 28924 22990 28926 23042
rect 28926 22990 28978 23042
rect 28978 22990 28980 23042
rect 28924 22988 28980 22990
rect 30380 23826 30436 23828
rect 30380 23774 30382 23826
rect 30382 23774 30434 23826
rect 30434 23774 30436 23826
rect 30380 23772 30436 23774
rect 27468 20242 27524 20244
rect 27468 20190 27470 20242
rect 27470 20190 27522 20242
rect 27522 20190 27524 20242
rect 27468 20188 27524 20190
rect 31164 20860 31220 20916
rect 29708 20188 29764 20244
rect 29820 20636 29876 20692
rect 30380 20690 30436 20692
rect 30380 20638 30382 20690
rect 30382 20638 30434 20690
rect 30434 20638 30436 20690
rect 30380 20636 30436 20638
rect 28812 19964 28868 20020
rect 30604 20076 30660 20132
rect 32172 23938 32228 23940
rect 32172 23886 32174 23938
rect 32174 23886 32226 23938
rect 32226 23886 32228 23938
rect 32172 23884 32228 23886
rect 31500 23826 31556 23828
rect 31500 23774 31502 23826
rect 31502 23774 31554 23826
rect 31554 23774 31556 23826
rect 31500 23772 31556 23774
rect 31836 23660 31892 23716
rect 32844 23714 32900 23716
rect 32844 23662 32846 23714
rect 32846 23662 32898 23714
rect 32898 23662 32900 23714
rect 32844 23660 32900 23662
rect 32396 23548 32452 23604
rect 32956 21644 33012 21700
rect 32508 20914 32564 20916
rect 32508 20862 32510 20914
rect 32510 20862 32562 20914
rect 32562 20862 32564 20914
rect 32508 20860 32564 20862
rect 32956 20188 33012 20244
rect 30940 20018 30996 20020
rect 30940 19966 30942 20018
rect 30942 19966 30994 20018
rect 30994 19966 30996 20018
rect 30940 19964 30996 19966
rect 36540 29314 36596 29316
rect 36540 29262 36542 29314
rect 36542 29262 36594 29314
rect 36594 29262 36596 29314
rect 36540 29260 36596 29262
rect 39116 29314 39172 29316
rect 39116 29262 39118 29314
rect 39118 29262 39170 29314
rect 39170 29262 39172 29314
rect 39116 29260 39172 29262
rect 38220 29148 38276 29204
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 34972 28754 35028 28756
rect 34972 28702 34974 28754
rect 34974 28702 35026 28754
rect 35026 28702 35028 28754
rect 34972 28700 35028 28702
rect 39228 29202 39284 29204
rect 39228 29150 39230 29202
rect 39230 29150 39282 29202
rect 39282 29150 39284 29202
rect 39228 29148 39284 29150
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35084 27074 35140 27076
rect 35084 27022 35086 27074
rect 35086 27022 35138 27074
rect 35138 27022 35140 27074
rect 35084 27020 35140 27022
rect 35756 27020 35812 27076
rect 34188 26684 34244 26740
rect 37884 27074 37940 27076
rect 37884 27022 37886 27074
rect 37886 27022 37938 27074
rect 37938 27022 37940 27074
rect 37884 27020 37940 27022
rect 41916 34130 41972 34132
rect 41916 34078 41918 34130
rect 41918 34078 41970 34130
rect 41970 34078 41972 34130
rect 41916 34076 41972 34078
rect 41580 33628 41636 33684
rect 42812 33628 42868 33684
rect 43596 35308 43652 35364
rect 46284 36540 46340 36596
rect 44716 35196 44772 35252
rect 44716 34914 44772 34916
rect 44716 34862 44718 34914
rect 44718 34862 44770 34914
rect 44770 34862 44772 34914
rect 44716 34860 44772 34862
rect 45276 34860 45332 34916
rect 45388 34018 45444 34020
rect 45388 33966 45390 34018
rect 45390 33966 45442 34018
rect 45442 33966 45444 34018
rect 45388 33964 45444 33966
rect 43820 32396 43876 32452
rect 44940 32396 44996 32452
rect 47628 39452 47684 39508
rect 49532 39452 49588 39508
rect 49868 39676 49924 39732
rect 49756 39116 49812 39172
rect 47740 38834 47796 38836
rect 47740 38782 47742 38834
rect 47742 38782 47794 38834
rect 47794 38782 47796 38834
rect 47740 38780 47796 38782
rect 48188 38668 48244 38724
rect 48188 38444 48244 38500
rect 48412 37212 48468 37268
rect 48748 38610 48804 38612
rect 48748 38558 48750 38610
rect 48750 38558 48802 38610
rect 48802 38558 48804 38610
rect 48748 38556 48804 38558
rect 49532 38834 49588 38836
rect 49532 38782 49534 38834
rect 49534 38782 49586 38834
rect 49586 38782 49588 38834
rect 49532 38780 49588 38782
rect 49756 38556 49812 38612
rect 48972 37212 49028 37268
rect 47852 37100 47908 37156
rect 46844 36540 46900 36596
rect 46956 36988 47012 37044
rect 48076 37042 48132 37044
rect 48076 36990 48078 37042
rect 48078 36990 48130 37042
rect 48130 36990 48132 37042
rect 48076 36988 48132 36990
rect 48412 37042 48468 37044
rect 48412 36990 48414 37042
rect 48414 36990 48466 37042
rect 48466 36990 48468 37042
rect 48412 36988 48468 36990
rect 49532 37266 49588 37268
rect 49532 37214 49534 37266
rect 49534 37214 49586 37266
rect 49586 37214 49588 37266
rect 49532 37212 49588 37214
rect 49756 37266 49812 37268
rect 49756 37214 49758 37266
rect 49758 37214 49810 37266
rect 49810 37214 49812 37266
rect 49756 37212 49812 37214
rect 54012 44322 54068 44324
rect 54012 44270 54014 44322
rect 54014 44270 54066 44322
rect 54066 44270 54068 44322
rect 54012 44268 54068 44270
rect 53004 43596 53060 43652
rect 53340 43596 53396 43652
rect 51884 42754 51940 42756
rect 51884 42702 51886 42754
rect 51886 42702 51938 42754
rect 51938 42702 51940 42754
rect 51884 42700 51940 42702
rect 53340 42194 53396 42196
rect 53340 42142 53342 42194
rect 53342 42142 53394 42194
rect 53394 42142 53396 42194
rect 53340 42140 53396 42142
rect 54124 42140 54180 42196
rect 51212 39618 51268 39620
rect 51212 39566 51214 39618
rect 51214 39566 51266 39618
rect 51266 39566 51268 39618
rect 51212 39564 51268 39566
rect 50092 39116 50148 39172
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 51212 39004 51268 39060
rect 49980 38444 50036 38500
rect 53676 39730 53732 39732
rect 53676 39678 53678 39730
rect 53678 39678 53730 39730
rect 53730 39678 53732 39730
rect 53676 39676 53732 39678
rect 52332 39564 52388 39620
rect 52332 38892 52388 38948
rect 51660 38834 51716 38836
rect 51660 38782 51662 38834
rect 51662 38782 51714 38834
rect 51714 38782 51716 38834
rect 51660 38780 51716 38782
rect 52444 38780 52500 38836
rect 50988 38668 51044 38724
rect 50652 38444 50708 38500
rect 51436 38722 51492 38724
rect 51436 38670 51438 38722
rect 51438 38670 51490 38722
rect 51490 38670 51492 38722
rect 51436 38668 51492 38670
rect 53676 39506 53732 39508
rect 53676 39454 53678 39506
rect 53678 39454 53730 39506
rect 53730 39454 53732 39506
rect 53676 39452 53732 39454
rect 53452 38892 53508 38948
rect 53004 38668 53060 38724
rect 53340 38722 53396 38724
rect 53340 38670 53342 38722
rect 53342 38670 53394 38722
rect 53394 38670 53396 38722
rect 53340 38668 53396 38670
rect 52108 38162 52164 38164
rect 52108 38110 52110 38162
rect 52110 38110 52162 38162
rect 52162 38110 52164 38162
rect 52108 38108 52164 38110
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 52892 38610 52948 38612
rect 52892 38558 52894 38610
rect 52894 38558 52946 38610
rect 52946 38558 52948 38610
rect 52892 38556 52948 38558
rect 52780 38108 52836 38164
rect 52556 37378 52612 37380
rect 52556 37326 52558 37378
rect 52558 37326 52610 37378
rect 52610 37326 52612 37378
rect 52556 37324 52612 37326
rect 51324 37266 51380 37268
rect 51324 37214 51326 37266
rect 51326 37214 51378 37266
rect 51378 37214 51380 37266
rect 51324 37212 51380 37214
rect 51548 37266 51604 37268
rect 51548 37214 51550 37266
rect 51550 37214 51602 37266
rect 51602 37214 51604 37266
rect 51548 37212 51604 37214
rect 52108 37154 52164 37156
rect 52108 37102 52110 37154
rect 52110 37102 52162 37154
rect 52162 37102 52164 37154
rect 52108 37100 52164 37102
rect 50092 36988 50148 37044
rect 54684 46508 54740 46564
rect 55132 44940 55188 44996
rect 55916 44994 55972 44996
rect 55916 44942 55918 44994
rect 55918 44942 55970 44994
rect 55970 44942 55972 44994
rect 55916 44940 55972 44942
rect 56252 43650 56308 43652
rect 56252 43598 56254 43650
rect 56254 43598 56306 43650
rect 56306 43598 56308 43650
rect 56252 43596 56308 43598
rect 54572 39676 54628 39732
rect 54012 38780 54068 38836
rect 54124 38722 54180 38724
rect 54124 38670 54126 38722
rect 54126 38670 54178 38722
rect 54178 38670 54180 38722
rect 54124 38668 54180 38670
rect 54236 38556 54292 38612
rect 54348 38108 54404 38164
rect 56364 38162 56420 38164
rect 56364 38110 56366 38162
rect 56366 38110 56418 38162
rect 56418 38110 56420 38162
rect 56364 38108 56420 38110
rect 53676 37378 53732 37380
rect 53676 37326 53678 37378
rect 53678 37326 53730 37378
rect 53730 37326 53732 37378
rect 53676 37324 53732 37326
rect 53564 37266 53620 37268
rect 53564 37214 53566 37266
rect 53566 37214 53618 37266
rect 53618 37214 53620 37266
rect 53564 37212 53620 37214
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 46844 34300 46900 34356
rect 47740 34354 47796 34356
rect 47740 34302 47742 34354
rect 47742 34302 47794 34354
rect 47794 34302 47796 34354
rect 47740 34300 47796 34302
rect 46284 33964 46340 34020
rect 48076 33964 48132 34020
rect 45612 32396 45668 32452
rect 46172 32450 46228 32452
rect 46172 32398 46174 32450
rect 46174 32398 46226 32450
rect 46226 32398 46228 32450
rect 46172 32396 46228 32398
rect 45388 31724 45444 31780
rect 44156 30210 44212 30212
rect 44156 30158 44158 30210
rect 44158 30158 44210 30210
rect 44210 30158 44212 30210
rect 44156 30156 44212 30158
rect 41580 29426 41636 29428
rect 41580 29374 41582 29426
rect 41582 29374 41634 29426
rect 41634 29374 41636 29426
rect 41580 29372 41636 29374
rect 45388 30156 45444 30212
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 46844 31778 46900 31780
rect 46844 31726 46846 31778
rect 46846 31726 46898 31778
rect 46898 31726 46900 31778
rect 46844 31724 46900 31726
rect 45948 30994 46004 30996
rect 45948 30942 45950 30994
rect 45950 30942 46002 30994
rect 46002 30942 46004 30994
rect 45948 30940 46004 30942
rect 48524 30322 48580 30324
rect 48524 30270 48526 30322
rect 48526 30270 48578 30322
rect 48578 30270 48580 30322
rect 48524 30268 48580 30270
rect 51212 31778 51268 31780
rect 51212 31726 51214 31778
rect 51214 31726 51266 31778
rect 51266 31726 51268 31778
rect 51212 31724 51268 31726
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 49532 30994 49588 30996
rect 49532 30942 49534 30994
rect 49534 30942 49586 30994
rect 49586 30942 49588 30994
rect 49532 30940 49588 30942
rect 49756 30434 49812 30436
rect 49756 30382 49758 30434
rect 49758 30382 49810 30434
rect 49810 30382 49812 30434
rect 49756 30380 49812 30382
rect 52444 30380 52500 30436
rect 49532 30322 49588 30324
rect 49532 30270 49534 30322
rect 49534 30270 49586 30322
rect 49586 30270 49588 30322
rect 49532 30268 49588 30270
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 41356 28700 41412 28756
rect 44492 29314 44548 29316
rect 44492 29262 44494 29314
rect 44494 29262 44546 29314
rect 44546 29262 44548 29314
rect 44492 29260 44548 29262
rect 45388 29314 45444 29316
rect 45388 29262 45390 29314
rect 45390 29262 45442 29314
rect 45442 29262 45444 29314
rect 45388 29260 45444 29262
rect 45948 29314 46004 29316
rect 45948 29262 45950 29314
rect 45950 29262 46002 29314
rect 46002 29262 46004 29314
rect 45948 29260 46004 29262
rect 49532 29314 49588 29316
rect 49532 29262 49534 29314
rect 49534 29262 49586 29314
rect 49586 29262 49588 29314
rect 49532 29260 49588 29262
rect 39788 27020 39844 27076
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 34748 25506 34804 25508
rect 34748 25454 34750 25506
rect 34750 25454 34802 25506
rect 34802 25454 34804 25506
rect 34748 25452 34804 25454
rect 34300 23938 34356 23940
rect 34300 23886 34302 23938
rect 34302 23886 34354 23938
rect 34354 23886 34356 23938
rect 34300 23884 34356 23886
rect 33628 23042 33684 23044
rect 33628 22990 33630 23042
rect 33630 22990 33682 23042
rect 33682 22990 33684 23042
rect 33628 22988 33684 22990
rect 33964 22652 34020 22708
rect 40236 26290 40292 26292
rect 40236 26238 40238 26290
rect 40238 26238 40290 26290
rect 40290 26238 40292 26290
rect 40236 26236 40292 26238
rect 40796 26124 40852 26180
rect 39788 26012 39844 26068
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34860 22988 34916 23044
rect 36204 23884 36260 23940
rect 36540 23884 36596 23940
rect 37548 23938 37604 23940
rect 37548 23886 37550 23938
rect 37550 23886 37602 23938
rect 37602 23886 37604 23938
rect 37548 23884 37604 23886
rect 38668 23660 38724 23716
rect 36764 23548 36820 23604
rect 34972 22652 35028 22708
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34636 22258 34692 22260
rect 34636 22206 34638 22258
rect 34638 22206 34690 22258
rect 34690 22206 34692 22258
rect 34636 22204 34692 22206
rect 33740 21644 33796 21700
rect 35756 22204 35812 22260
rect 35084 21644 35140 21700
rect 35644 21698 35700 21700
rect 35644 21646 35646 21698
rect 35646 21646 35698 21698
rect 35698 21646 35700 21698
rect 35644 21644 35700 21646
rect 34972 21586 35028 21588
rect 34972 21534 34974 21586
rect 34974 21534 35026 21586
rect 35026 21534 35028 21586
rect 34972 21532 35028 21534
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 33964 20188 34020 20244
rect 35644 20524 35700 20580
rect 34860 20188 34916 20244
rect 33404 18396 33460 18452
rect 27580 17106 27636 17108
rect 27580 17054 27582 17106
rect 27582 17054 27634 17106
rect 27634 17054 27636 17106
rect 27580 17052 27636 17054
rect 28140 17052 28196 17108
rect 27916 14588 27972 14644
rect 26236 13468 26292 13524
rect 36540 20076 36596 20132
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 33516 18284 33572 18340
rect 34636 18284 34692 18340
rect 29036 17052 29092 17108
rect 31052 16828 31108 16884
rect 32956 16940 33012 16996
rect 33740 16994 33796 16996
rect 33740 16942 33742 16994
rect 33742 16942 33794 16994
rect 33794 16942 33796 16994
rect 33740 16940 33796 16942
rect 33628 16882 33684 16884
rect 33628 16830 33630 16882
rect 33630 16830 33682 16882
rect 33682 16830 33684 16882
rect 33628 16828 33684 16830
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34748 17106 34804 17108
rect 34748 17054 34750 17106
rect 34750 17054 34802 17106
rect 34802 17054 34804 17106
rect 34748 17052 34804 17054
rect 43484 27858 43540 27860
rect 43484 27806 43486 27858
rect 43486 27806 43538 27858
rect 43538 27806 43540 27858
rect 43484 27804 43540 27806
rect 46508 27804 46564 27860
rect 41804 27074 41860 27076
rect 41804 27022 41806 27074
rect 41806 27022 41858 27074
rect 41858 27022 41860 27074
rect 41804 27020 41860 27022
rect 46732 27858 46788 27860
rect 46732 27806 46734 27858
rect 46734 27806 46786 27858
rect 46786 27806 46788 27858
rect 46732 27804 46788 27806
rect 48076 27858 48132 27860
rect 48076 27806 48078 27858
rect 48078 27806 48130 27858
rect 48130 27806 48132 27858
rect 48076 27804 48132 27806
rect 40124 25506 40180 25508
rect 40124 25454 40126 25506
rect 40126 25454 40178 25506
rect 40178 25454 40180 25506
rect 40124 25452 40180 25454
rect 41020 23714 41076 23716
rect 41020 23662 41022 23714
rect 41022 23662 41074 23714
rect 41074 23662 41076 23714
rect 41020 23660 41076 23662
rect 37996 22370 38052 22372
rect 37996 22318 37998 22370
rect 37998 22318 38050 22370
rect 38050 22318 38052 22370
rect 37996 22316 38052 22318
rect 39228 22316 39284 22372
rect 42364 26460 42420 26516
rect 48524 26908 48580 26964
rect 42028 26178 42084 26180
rect 42028 26126 42030 26178
rect 42030 26126 42082 26178
rect 42082 26126 42084 26178
rect 42028 26124 42084 26126
rect 41804 26066 41860 26068
rect 41804 26014 41806 26066
rect 41806 26014 41858 26066
rect 41858 26014 41860 26066
rect 41804 26012 41860 26014
rect 42812 26236 42868 26292
rect 41804 25452 41860 25508
rect 41804 24780 41860 24836
rect 42588 24556 42644 24612
rect 42028 23154 42084 23156
rect 42028 23102 42030 23154
rect 42030 23102 42082 23154
rect 42082 23102 42084 23154
rect 42028 23100 42084 23102
rect 39228 21644 39284 21700
rect 41468 21698 41524 21700
rect 41468 21646 41470 21698
rect 41470 21646 41522 21698
rect 41522 21646 41524 21698
rect 41468 21644 41524 21646
rect 39340 21586 39396 21588
rect 39340 21534 39342 21586
rect 39342 21534 39394 21586
rect 39394 21534 39396 21586
rect 39340 21532 39396 21534
rect 37548 20578 37604 20580
rect 37548 20526 37550 20578
rect 37550 20526 37602 20578
rect 37602 20526 37604 20578
rect 37548 20524 37604 20526
rect 37436 20188 37492 20244
rect 36988 19964 37044 20020
rect 38108 20188 38164 20244
rect 38444 20130 38500 20132
rect 38444 20078 38446 20130
rect 38446 20078 38498 20130
rect 38498 20078 38500 20130
rect 38444 20076 38500 20078
rect 38332 20018 38388 20020
rect 38332 19966 38334 20018
rect 38334 19966 38386 20018
rect 38386 19966 38388 20018
rect 38332 19964 38388 19966
rect 37772 19906 37828 19908
rect 37772 19854 37774 19906
rect 37774 19854 37826 19906
rect 37826 19854 37828 19906
rect 37772 19852 37828 19854
rect 38108 19234 38164 19236
rect 38108 19182 38110 19234
rect 38110 19182 38162 19234
rect 38162 19182 38164 19234
rect 38108 19180 38164 19182
rect 40012 20188 40068 20244
rect 40572 20242 40628 20244
rect 40572 20190 40574 20242
rect 40574 20190 40626 20242
rect 40626 20190 40628 20242
rect 40572 20188 40628 20190
rect 39340 19852 39396 19908
rect 44716 25394 44772 25396
rect 44716 25342 44718 25394
rect 44718 25342 44770 25394
rect 44770 25342 44772 25394
rect 44716 25340 44772 25342
rect 45500 25394 45556 25396
rect 45500 25342 45502 25394
rect 45502 25342 45554 25394
rect 45554 25342 45556 25394
rect 45500 25340 45556 25342
rect 44492 25282 44548 25284
rect 44492 25230 44494 25282
rect 44494 25230 44546 25282
rect 44546 25230 44548 25282
rect 44492 25228 44548 25230
rect 45388 25228 45444 25284
rect 43708 24892 43764 24948
rect 44940 24946 44996 24948
rect 44940 24894 44942 24946
rect 44942 24894 44994 24946
rect 44994 24894 44996 24946
rect 44940 24892 44996 24894
rect 44716 24050 44772 24052
rect 44716 23998 44718 24050
rect 44718 23998 44770 24050
rect 44770 23998 44772 24050
rect 44716 23996 44772 23998
rect 45612 24610 45668 24612
rect 45612 24558 45614 24610
rect 45614 24558 45666 24610
rect 45666 24558 45668 24610
rect 45612 24556 45668 24558
rect 42812 23100 42868 23156
rect 42028 21532 42084 21588
rect 42140 21644 42196 21700
rect 43484 21532 43540 21588
rect 42924 21474 42980 21476
rect 42924 21422 42926 21474
rect 42926 21422 42978 21474
rect 42978 21422 42980 21474
rect 42924 21420 42980 21422
rect 41468 20076 41524 20132
rect 39900 19292 39956 19348
rect 40908 19346 40964 19348
rect 40908 19294 40910 19346
rect 40910 19294 40962 19346
rect 40962 19294 40964 19346
rect 40908 19292 40964 19294
rect 45052 21474 45108 21476
rect 45052 21422 45054 21474
rect 45054 21422 45106 21474
rect 45106 21422 45108 21474
rect 45052 21420 45108 21422
rect 45612 22316 45668 22372
rect 47516 26178 47572 26180
rect 47516 26126 47518 26178
rect 47518 26126 47570 26178
rect 47570 26126 47572 26178
rect 47516 26124 47572 26126
rect 48860 26348 48916 26404
rect 48748 26290 48804 26292
rect 48748 26238 48750 26290
rect 48750 26238 48802 26290
rect 48802 26238 48804 26290
rect 48748 26236 48804 26238
rect 48748 25506 48804 25508
rect 48748 25454 48750 25506
rect 48750 25454 48802 25506
rect 48802 25454 48804 25506
rect 48748 25452 48804 25454
rect 48076 25228 48132 25284
rect 48412 25282 48468 25284
rect 48412 25230 48414 25282
rect 48414 25230 48466 25282
rect 48466 25230 48468 25282
rect 48412 25228 48468 25230
rect 46844 24892 46900 24948
rect 47068 23996 47124 24052
rect 46396 23548 46452 23604
rect 46620 23324 46676 23380
rect 45836 22204 45892 22260
rect 45612 21420 45668 21476
rect 45164 20748 45220 20804
rect 42588 20076 42644 20132
rect 41356 19180 41412 19236
rect 28476 13186 28532 13188
rect 28476 13134 28478 13186
rect 28478 13134 28530 13186
rect 28530 13134 28532 13186
rect 28476 13132 28532 13134
rect 29036 13132 29092 13188
rect 29148 13468 29204 13524
rect 26124 11564 26180 11620
rect 28028 12178 28084 12180
rect 28028 12126 28030 12178
rect 28030 12126 28082 12178
rect 28082 12126 28084 12178
rect 28028 12124 28084 12126
rect 26348 11452 26404 11508
rect 28364 11954 28420 11956
rect 28364 11902 28366 11954
rect 28366 11902 28418 11954
rect 28418 11902 28420 11954
rect 28364 11900 28420 11902
rect 32060 13916 32116 13972
rect 29820 11788 29876 11844
rect 26908 9266 26964 9268
rect 26908 9214 26910 9266
rect 26910 9214 26962 9266
rect 26962 9214 26964 9266
rect 26908 9212 26964 9214
rect 27580 9826 27636 9828
rect 27580 9774 27582 9826
rect 27582 9774 27634 9826
rect 27634 9774 27636 9826
rect 27580 9772 27636 9774
rect 33516 13970 33572 13972
rect 33516 13918 33518 13970
rect 33518 13918 33570 13970
rect 33570 13918 33572 13970
rect 33516 13916 33572 13918
rect 37324 17052 37380 17108
rect 36764 16828 36820 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 40796 18450 40852 18452
rect 40796 18398 40798 18450
rect 40798 18398 40850 18450
rect 40850 18398 40852 18450
rect 40796 18396 40852 18398
rect 41916 18450 41972 18452
rect 41916 18398 41918 18450
rect 41918 18398 41970 18450
rect 41970 18398 41972 18450
rect 41916 18396 41972 18398
rect 41020 17554 41076 17556
rect 41020 17502 41022 17554
rect 41022 17502 41074 17554
rect 41074 17502 41076 17554
rect 41020 17500 41076 17502
rect 38556 16882 38612 16884
rect 38556 16830 38558 16882
rect 38558 16830 38610 16882
rect 38610 16830 38612 16882
rect 38556 16828 38612 16830
rect 37772 16210 37828 16212
rect 37772 16158 37774 16210
rect 37774 16158 37826 16210
rect 37826 16158 37828 16210
rect 37772 16156 37828 16158
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 34076 13916 34132 13972
rect 35308 13916 35364 13972
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 31948 11788 32004 11844
rect 32172 11900 32228 11956
rect 35644 12908 35700 12964
rect 36316 12962 36372 12964
rect 36316 12910 36318 12962
rect 36318 12910 36370 12962
rect 36370 12910 36372 12962
rect 36316 12908 36372 12910
rect 33964 12402 34020 12404
rect 33964 12350 33966 12402
rect 33966 12350 34018 12402
rect 34018 12350 34020 12402
rect 33964 12348 34020 12350
rect 35532 12348 35588 12404
rect 36988 12348 37044 12404
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 38332 11618 38388 11620
rect 38332 11566 38334 11618
rect 38334 11566 38386 11618
rect 38386 11566 38388 11618
rect 38332 11564 38388 11566
rect 35756 11452 35812 11508
rect 36204 11506 36260 11508
rect 36204 11454 36206 11506
rect 36206 11454 36258 11506
rect 36258 11454 36260 11506
rect 36204 11452 36260 11454
rect 38780 16210 38836 16212
rect 38780 16158 38782 16210
rect 38782 16158 38834 16210
rect 38834 16158 38836 16210
rect 38780 16156 38836 16158
rect 39788 16156 39844 16212
rect 40908 16210 40964 16212
rect 40908 16158 40910 16210
rect 40910 16158 40962 16210
rect 40962 16158 40964 16210
rect 40908 16156 40964 16158
rect 42364 17554 42420 17556
rect 42364 17502 42366 17554
rect 42366 17502 42418 17554
rect 42418 17502 42420 17554
rect 42364 17500 42420 17502
rect 43932 20076 43988 20132
rect 46284 22316 46340 22372
rect 46508 22258 46564 22260
rect 46508 22206 46510 22258
rect 46510 22206 46562 22258
rect 46562 22206 46564 22258
rect 46508 22204 46564 22206
rect 46060 21868 46116 21924
rect 45948 20802 46004 20804
rect 45948 20750 45950 20802
rect 45950 20750 46002 20802
rect 46002 20750 46004 20802
rect 45948 20748 46004 20750
rect 47964 23660 48020 23716
rect 47740 23436 47796 23492
rect 47180 22594 47236 22596
rect 47180 22542 47182 22594
rect 47182 22542 47234 22594
rect 47234 22542 47236 22594
rect 47180 22540 47236 22542
rect 47068 22316 47124 22372
rect 47404 22652 47460 22708
rect 47180 21868 47236 21924
rect 48076 23324 48132 23380
rect 48076 22652 48132 22708
rect 49756 27804 49812 27860
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 49756 26908 49812 26964
rect 49644 26348 49700 26404
rect 49532 26290 49588 26292
rect 49532 26238 49534 26290
rect 49534 26238 49586 26290
rect 49586 26238 49588 26290
rect 49532 26236 49588 26238
rect 49868 26402 49924 26404
rect 49868 26350 49870 26402
rect 49870 26350 49922 26402
rect 49922 26350 49924 26402
rect 49868 26348 49924 26350
rect 49644 25564 49700 25620
rect 49868 25452 49924 25508
rect 49532 25394 49588 25396
rect 49532 25342 49534 25394
rect 49534 25342 49586 25394
rect 49586 25342 49588 25394
rect 49532 25340 49588 25342
rect 49532 23660 49588 23716
rect 48300 23100 48356 23156
rect 48300 22540 48356 22596
rect 47964 22370 48020 22372
rect 47964 22318 47966 22370
rect 47966 22318 48018 22370
rect 48018 22318 48020 22370
rect 47964 22316 48020 22318
rect 48076 21980 48132 22036
rect 47628 21532 47684 21588
rect 47180 20076 47236 20132
rect 42812 16882 42868 16884
rect 42812 16830 42814 16882
rect 42814 16830 42866 16882
rect 42866 16830 42868 16882
rect 42812 16828 42868 16830
rect 38892 15820 38948 15876
rect 44044 15986 44100 15988
rect 44044 15934 44046 15986
rect 44046 15934 44098 15986
rect 44098 15934 44100 15986
rect 44044 15932 44100 15934
rect 41692 15820 41748 15876
rect 39564 14588 39620 14644
rect 42140 15874 42196 15876
rect 42140 15822 42142 15874
rect 42142 15822 42194 15874
rect 42194 15822 42196 15874
rect 42140 15820 42196 15822
rect 39116 12962 39172 12964
rect 39116 12910 39118 12962
rect 39118 12910 39170 12962
rect 39170 12910 39172 12962
rect 39116 12908 39172 12910
rect 38892 12348 38948 12404
rect 38556 11564 38612 11620
rect 39116 11564 39172 11620
rect 41916 13074 41972 13076
rect 41916 13022 41918 13074
rect 41918 13022 41970 13074
rect 41970 13022 41972 13074
rect 41916 13020 41972 13022
rect 41580 12908 41636 12964
rect 40236 12402 40292 12404
rect 40236 12350 40238 12402
rect 40238 12350 40290 12402
rect 40290 12350 40292 12402
rect 40236 12348 40292 12350
rect 45388 16828 45444 16884
rect 46060 16882 46116 16884
rect 46060 16830 46062 16882
rect 46062 16830 46114 16882
rect 46114 16830 46116 16882
rect 46060 16828 46116 16830
rect 44716 15874 44772 15876
rect 44716 15822 44718 15874
rect 44718 15822 44770 15874
rect 44770 15822 44772 15874
rect 44716 15820 44772 15822
rect 44492 15260 44548 15316
rect 45612 15314 45668 15316
rect 45612 15262 45614 15314
rect 45614 15262 45666 15314
rect 45666 15262 45668 15314
rect 45612 15260 45668 15262
rect 46508 17724 46564 17780
rect 50204 26684 50260 26740
rect 50652 26850 50708 26852
rect 50652 26798 50654 26850
rect 50654 26798 50706 26850
rect 50706 26798 50708 26850
rect 50652 26796 50708 26798
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50428 25618 50484 25620
rect 50428 25566 50430 25618
rect 50430 25566 50482 25618
rect 50482 25566 50484 25618
rect 50428 25564 50484 25566
rect 50988 26348 51044 26404
rect 50876 25394 50932 25396
rect 50876 25342 50878 25394
rect 50878 25342 50930 25394
rect 50930 25342 50932 25394
rect 50876 25340 50932 25342
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 51100 26236 51156 26292
rect 52108 27804 52164 27860
rect 53340 27804 53396 27860
rect 51660 27074 51716 27076
rect 51660 27022 51662 27074
rect 51662 27022 51714 27074
rect 51714 27022 51716 27074
rect 51660 27020 51716 27022
rect 51548 26962 51604 26964
rect 51548 26910 51550 26962
rect 51550 26910 51602 26962
rect 51602 26910 51604 26962
rect 51548 26908 51604 26910
rect 52332 26962 52388 26964
rect 52332 26910 52334 26962
rect 52334 26910 52386 26962
rect 52386 26910 52388 26962
rect 52332 26908 52388 26910
rect 51324 26402 51380 26404
rect 51324 26350 51326 26402
rect 51326 26350 51378 26402
rect 51378 26350 51380 26402
rect 51324 26348 51380 26350
rect 51436 26290 51492 26292
rect 51436 26238 51438 26290
rect 51438 26238 51490 26290
rect 51490 26238 51492 26290
rect 51436 26236 51492 26238
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 49756 23154 49812 23156
rect 49756 23102 49758 23154
rect 49758 23102 49810 23154
rect 49810 23102 49812 23154
rect 49756 23100 49812 23102
rect 49644 21868 49700 21924
rect 51212 24722 51268 24724
rect 51212 24670 51214 24722
rect 51214 24670 51266 24722
rect 51266 24670 51268 24722
rect 51212 24668 51268 24670
rect 51548 24668 51604 24724
rect 53676 26796 53732 26852
rect 55356 26908 55412 26964
rect 52444 24668 52500 24724
rect 52668 24162 52724 24164
rect 52668 24110 52670 24162
rect 52670 24110 52722 24162
rect 52722 24110 52724 24162
rect 52668 24108 52724 24110
rect 54572 24108 54628 24164
rect 55356 24556 55412 24612
rect 50988 23100 51044 23156
rect 51100 23324 51156 23380
rect 50428 22876 50484 22932
rect 51100 22316 51156 22372
rect 51660 23660 51716 23716
rect 51548 22930 51604 22932
rect 51548 22878 51550 22930
rect 51550 22878 51602 22930
rect 51602 22878 51604 22930
rect 51548 22876 51604 22878
rect 52556 23714 52612 23716
rect 52556 23662 52558 23714
rect 52558 23662 52610 23714
rect 52610 23662 52612 23714
rect 52556 23660 52612 23662
rect 52220 23324 52276 23380
rect 51772 23100 51828 23156
rect 51436 22370 51492 22372
rect 51436 22318 51438 22370
rect 51438 22318 51490 22370
rect 51490 22318 51492 22370
rect 51436 22316 51492 22318
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50876 21810 50932 21812
rect 50876 21758 50878 21810
rect 50878 21758 50930 21810
rect 50930 21758 50932 21810
rect 50876 21756 50932 21758
rect 51436 21756 51492 21812
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 49644 20188 49700 20244
rect 50540 20242 50596 20244
rect 50540 20190 50542 20242
rect 50542 20190 50594 20242
rect 50594 20190 50596 20242
rect 50540 20188 50596 20190
rect 47628 17778 47684 17780
rect 47628 17726 47630 17778
rect 47630 17726 47682 17778
rect 47682 17726 47684 17778
rect 47628 17724 47684 17726
rect 47180 17052 47236 17108
rect 43820 14642 43876 14644
rect 43820 14590 43822 14642
rect 43822 14590 43874 14642
rect 43874 14590 43876 14642
rect 43820 14588 43876 14590
rect 45836 13020 45892 13076
rect 44044 12850 44100 12852
rect 44044 12798 44046 12850
rect 44046 12798 44098 12850
rect 44098 12798 44100 12850
rect 44044 12796 44100 12798
rect 41580 12178 41636 12180
rect 41580 12126 41582 12178
rect 41582 12126 41634 12178
rect 41634 12126 41636 12178
rect 41580 12124 41636 12126
rect 39564 11452 39620 11508
rect 45276 12124 45332 12180
rect 38556 11170 38612 11172
rect 38556 11118 38558 11170
rect 38558 11118 38610 11170
rect 38610 11118 38612 11170
rect 38556 11116 38612 11118
rect 39228 11116 39284 11172
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 39788 11116 39844 11172
rect 40012 11564 40068 11620
rect 44492 11564 44548 11620
rect 45724 11618 45780 11620
rect 45724 11566 45726 11618
rect 45726 11566 45778 11618
rect 45778 11566 45780 11618
rect 45724 11564 45780 11566
rect 46284 13020 46340 13076
rect 46284 12850 46340 12852
rect 46284 12798 46286 12850
rect 46286 12798 46338 12850
rect 46338 12798 46340 12850
rect 46284 12796 46340 12798
rect 46396 12348 46452 12404
rect 46060 11788 46116 11844
rect 46396 11788 46452 11844
rect 48300 17388 48356 17444
rect 48860 17442 48916 17444
rect 48860 17390 48862 17442
rect 48862 17390 48914 17442
rect 48914 17390 48916 17442
rect 48860 17388 48916 17390
rect 49644 18450 49700 18452
rect 49644 18398 49646 18450
rect 49646 18398 49698 18450
rect 49698 18398 49700 18450
rect 49644 18396 49700 18398
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 52780 23154 52836 23156
rect 52780 23102 52782 23154
rect 52782 23102 52834 23154
rect 52834 23102 52836 23154
rect 52780 23100 52836 23102
rect 52556 22876 52612 22932
rect 55916 24610 55972 24612
rect 55916 24558 55918 24610
rect 55918 24558 55970 24610
rect 55970 24558 55972 24610
rect 55916 24556 55972 24558
rect 51996 21196 52052 21252
rect 53676 21196 53732 21252
rect 51324 18396 51380 18452
rect 49644 17388 49700 17444
rect 48748 17106 48804 17108
rect 48748 17054 48750 17106
rect 48750 17054 48802 17106
rect 48802 17054 48804 17106
rect 48748 17052 48804 17054
rect 49532 17052 49588 17108
rect 47628 15986 47684 15988
rect 47628 15934 47630 15986
rect 47630 15934 47682 15986
rect 47682 15934 47684 15986
rect 47628 15932 47684 15934
rect 52668 19122 52724 19124
rect 52668 19070 52670 19122
rect 52670 19070 52722 19122
rect 52722 19070 52724 19122
rect 52668 19068 52724 19070
rect 54908 19180 54964 19236
rect 56252 19234 56308 19236
rect 56252 19182 56254 19234
rect 56254 19182 56306 19234
rect 56306 19182 56308 19234
rect 56252 19180 56308 19182
rect 56812 19234 56868 19236
rect 56812 19182 56814 19234
rect 56814 19182 56866 19234
rect 56866 19182 56868 19234
rect 56812 19180 56868 19182
rect 55580 19122 55636 19124
rect 55580 19070 55582 19122
rect 55582 19070 55634 19122
rect 55634 19070 55636 19122
rect 55580 19068 55636 19070
rect 51772 18172 51828 18228
rect 53228 18226 53284 18228
rect 53228 18174 53230 18226
rect 53230 18174 53282 18226
rect 53282 18174 53284 18226
rect 53228 18172 53284 18174
rect 51996 17442 52052 17444
rect 51996 17390 51998 17442
rect 51998 17390 52050 17442
rect 52050 17390 52052 17442
rect 51996 17388 52052 17390
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 52668 17442 52724 17444
rect 52668 17390 52670 17442
rect 52670 17390 52722 17442
rect 52722 17390 52724 17442
rect 52668 17388 52724 17390
rect 46956 14588 47012 14644
rect 49196 15372 49252 15428
rect 50540 15986 50596 15988
rect 50540 15934 50542 15986
rect 50542 15934 50594 15986
rect 50594 15934 50596 15986
rect 50540 15932 50596 15934
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50316 15426 50372 15428
rect 50316 15374 50318 15426
rect 50318 15374 50370 15426
rect 50370 15374 50372 15426
rect 50316 15372 50372 15374
rect 50316 14642 50372 14644
rect 50316 14590 50318 14642
rect 50318 14590 50370 14642
rect 50370 14590 50372 14642
rect 50316 14588 50372 14590
rect 46956 13746 47012 13748
rect 46956 13694 46958 13746
rect 46958 13694 47010 13746
rect 47010 13694 47012 13746
rect 46956 13692 47012 13694
rect 47852 13746 47908 13748
rect 47852 13694 47854 13746
rect 47854 13694 47906 13746
rect 47906 13694 47908 13746
rect 47852 13692 47908 13694
rect 47628 13020 47684 13076
rect 47516 11394 47572 11396
rect 47516 11342 47518 11394
rect 47518 11342 47570 11394
rect 47570 11342 47572 11394
rect 47516 11340 47572 11342
rect 46396 11282 46452 11284
rect 46396 11230 46398 11282
rect 46398 11230 46450 11282
rect 46450 11230 46452 11282
rect 46396 11228 46452 11230
rect 47404 11282 47460 11284
rect 47404 11230 47406 11282
rect 47406 11230 47458 11282
rect 47458 11230 47460 11282
rect 47404 11228 47460 11230
rect 45948 11116 46004 11172
rect 31948 9884 32004 9940
rect 38332 10108 38388 10164
rect 33068 9938 33124 9940
rect 33068 9886 33070 9938
rect 33070 9886 33122 9938
rect 33122 9886 33124 9938
rect 33068 9884 33124 9886
rect 24444 8204 24500 8260
rect 24668 7586 24724 7588
rect 24668 7534 24670 7586
rect 24670 7534 24722 7586
rect 24722 7534 24724 7586
rect 24668 7532 24724 7534
rect 24444 7250 24500 7252
rect 24444 7198 24446 7250
rect 24446 7198 24498 7250
rect 24498 7198 24500 7250
rect 24444 7196 24500 7198
rect 25564 7196 25620 7252
rect 26236 7586 26292 7588
rect 26236 7534 26238 7586
rect 26238 7534 26290 7586
rect 26290 7534 26292 7586
rect 26236 7532 26292 7534
rect 26572 7474 26628 7476
rect 26572 7422 26574 7474
rect 26574 7422 26626 7474
rect 26626 7422 26628 7474
rect 26572 7420 26628 7422
rect 27132 7420 27188 7476
rect 26796 7196 26852 7252
rect 27356 7196 27412 7252
rect 27804 7532 27860 7588
rect 37660 8988 37716 9044
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 27916 7420 27972 7476
rect 29932 7644 29988 7700
rect 30492 7698 30548 7700
rect 30492 7646 30494 7698
rect 30494 7646 30546 7698
rect 30546 7646 30548 7698
rect 30492 7644 30548 7646
rect 27804 7308 27860 7364
rect 26572 6636 26628 6692
rect 27244 6690 27300 6692
rect 27244 6638 27246 6690
rect 27246 6638 27298 6690
rect 27298 6638 27300 6690
rect 27244 6636 27300 6638
rect 29260 7362 29316 7364
rect 29260 7310 29262 7362
rect 29262 7310 29314 7362
rect 29314 7310 29316 7362
rect 29260 7308 29316 7310
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 38780 10108 38836 10164
rect 38220 7474 38276 7476
rect 38220 7422 38222 7474
rect 38222 7422 38274 7474
rect 38274 7422 38276 7474
rect 38220 7420 38276 7422
rect 38780 7420 38836 7476
rect 39228 7420 39284 7476
rect 38556 7362 38612 7364
rect 38556 7310 38558 7362
rect 38558 7310 38610 7362
rect 38610 7310 38612 7362
rect 38556 7308 38612 7310
rect 39116 7362 39172 7364
rect 39116 7310 39118 7362
rect 39118 7310 39170 7362
rect 39170 7310 39172 7362
rect 39116 7308 39172 7310
rect 23660 6076 23716 6132
rect 26236 6130 26292 6132
rect 26236 6078 26238 6130
rect 26238 6078 26290 6130
rect 26290 6078 26292 6130
rect 26236 6076 26292 6078
rect 39564 9884 39620 9940
rect 40460 9938 40516 9940
rect 40460 9886 40462 9938
rect 40462 9886 40514 9938
rect 40514 9886 40516 9938
rect 40460 9884 40516 9886
rect 40236 9042 40292 9044
rect 40236 8990 40238 9042
rect 40238 8990 40290 9042
rect 40290 8990 40292 9042
rect 40236 8988 40292 8990
rect 40684 9042 40740 9044
rect 40684 8990 40686 9042
rect 40686 8990 40738 9042
rect 40738 8990 40740 9042
rect 40684 8988 40740 8990
rect 47180 11170 47236 11172
rect 47180 11118 47182 11170
rect 47182 11118 47234 11170
rect 47234 11118 47236 11170
rect 47180 11116 47236 11118
rect 44716 10332 44772 10388
rect 41020 8988 41076 9044
rect 41804 9042 41860 9044
rect 41804 8990 41806 9042
rect 41806 8990 41858 9042
rect 41858 8990 41860 9042
rect 41804 8988 41860 8990
rect 44380 8876 44436 8932
rect 44604 9212 44660 9268
rect 45388 10386 45444 10388
rect 45388 10334 45390 10386
rect 45390 10334 45442 10386
rect 45442 10334 45444 10386
rect 45388 10332 45444 10334
rect 45164 9996 45220 10052
rect 45164 9266 45220 9268
rect 45164 9214 45166 9266
rect 45166 9214 45218 9266
rect 45218 9214 45220 9266
rect 45164 9212 45220 9214
rect 43260 7586 43316 7588
rect 43260 7534 43262 7586
rect 43262 7534 43314 7586
rect 43314 7534 43316 7586
rect 43260 7532 43316 7534
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 53452 15986 53508 15988
rect 53452 15934 53454 15986
rect 53454 15934 53506 15986
rect 53506 15934 53508 15986
rect 53452 15932 53508 15934
rect 54796 17724 54852 17780
rect 55916 17778 55972 17780
rect 55916 17726 55918 17778
rect 55918 17726 55970 17778
rect 55970 17726 55972 17778
rect 55916 17724 55972 17726
rect 52780 13692 52836 13748
rect 53116 14588 53172 14644
rect 53564 13746 53620 13748
rect 53564 13694 53566 13746
rect 53566 13694 53618 13746
rect 53618 13694 53620 13746
rect 53564 13692 53620 13694
rect 54124 14588 54180 14644
rect 55580 14642 55636 14644
rect 55580 14590 55582 14642
rect 55582 14590 55634 14642
rect 55634 14590 55636 14642
rect 55580 14588 55636 14590
rect 48412 12348 48468 12404
rect 52220 12684 52276 12740
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50764 11564 50820 11620
rect 51996 11676 52052 11732
rect 50988 11506 51044 11508
rect 50988 11454 50990 11506
rect 50990 11454 51042 11506
rect 51042 11454 51044 11506
rect 50988 11452 51044 11454
rect 47852 9996 47908 10052
rect 48076 9996 48132 10052
rect 46620 9884 46676 9940
rect 47628 9938 47684 9940
rect 47628 9886 47630 9938
rect 47630 9886 47682 9938
rect 47682 9886 47684 9938
rect 47628 9884 47684 9886
rect 51996 11394 52052 11396
rect 51996 11342 51998 11394
rect 51998 11342 52050 11394
rect 52050 11342 52052 11394
rect 51996 11340 52052 11342
rect 53340 12738 53396 12740
rect 53340 12686 53342 12738
rect 53342 12686 53394 12738
rect 53394 12686 53396 12738
rect 53340 12684 53396 12686
rect 53676 12348 53732 12404
rect 53564 11618 53620 11620
rect 53564 11566 53566 11618
rect 53566 11566 53618 11618
rect 53618 11566 53620 11618
rect 53564 11564 53620 11566
rect 53676 11506 53732 11508
rect 53676 11454 53678 11506
rect 53678 11454 53730 11506
rect 53730 11454 53732 11506
rect 53676 11452 53732 11454
rect 53452 11340 53508 11396
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50876 10556 50932 10612
rect 51436 10610 51492 10612
rect 51436 10558 51438 10610
rect 51438 10558 51490 10610
rect 51490 10558 51492 10610
rect 51436 10556 51492 10558
rect 50876 9996 50932 10052
rect 48636 9548 48692 9604
rect 50316 9548 50372 9604
rect 48748 8204 48804 8260
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 52444 10108 52500 10164
rect 53900 10108 53956 10164
rect 49084 8316 49140 8372
rect 54460 12684 54516 12740
rect 55020 12402 55076 12404
rect 55020 12350 55022 12402
rect 55022 12350 55074 12402
rect 55074 12350 55076 12402
rect 55020 12348 55076 12350
rect 56364 12348 56420 12404
rect 54236 11788 54292 11844
rect 54124 11394 54180 11396
rect 54124 11342 54126 11394
rect 54126 11342 54178 11394
rect 54178 11342 54180 11394
rect 54124 11340 54180 11342
rect 51324 8316 51380 8372
rect 51772 8316 51828 8372
rect 45500 7532 45556 7588
rect 39788 6636 39844 6692
rect 40012 6636 40068 6692
rect 40460 6636 40516 6692
rect 28 3612 84 3668
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 2492 3666 2548 3668
rect 2492 3614 2494 3666
rect 2494 3614 2546 3666
rect 2546 3614 2548 3666
rect 2492 3612 2548 3614
rect 21532 3612 21588 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 40124 5180 40180 5236
rect 40572 5122 40628 5124
rect 40572 5070 40574 5122
rect 40574 5070 40626 5122
rect 40626 5070 40628 5122
rect 40572 5068 40628 5070
rect 41244 5234 41300 5236
rect 41244 5182 41246 5234
rect 41246 5182 41298 5234
rect 41298 5182 41300 5234
rect 41244 5180 41300 5182
rect 40908 5068 40964 5124
rect 46284 6748 46340 6804
rect 49756 8258 49812 8260
rect 49756 8206 49758 8258
rect 49758 8206 49810 8258
rect 49810 8206 49812 8258
rect 49756 8204 49812 8206
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 51884 8204 51940 8260
rect 52668 8370 52724 8372
rect 52668 8318 52670 8370
rect 52670 8318 52722 8370
rect 52722 8318 52724 8370
rect 52668 8316 52724 8318
rect 48972 6748 49028 6804
rect 49084 6636 49140 6692
rect 49420 6748 49476 6804
rect 49644 6748 49700 6804
rect 52332 7362 52388 7364
rect 52332 7310 52334 7362
rect 52334 7310 52386 7362
rect 52386 7310 52388 7362
rect 52332 7308 52388 7310
rect 52556 6860 52612 6916
rect 53564 7308 53620 7364
rect 53788 6860 53844 6916
rect 52668 6748 52724 6804
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 53340 6802 53396 6804
rect 53340 6750 53342 6802
rect 53342 6750 53394 6802
rect 53394 6750 53396 6802
rect 53340 6748 53396 6750
rect 54124 8258 54180 8260
rect 54124 8206 54126 8258
rect 54126 8206 54178 8258
rect 54178 8206 54180 8258
rect 54124 8204 54180 8206
rect 54460 7586 54516 7588
rect 54460 7534 54462 7586
rect 54462 7534 54514 7586
rect 54514 7534 54516 7586
rect 54460 7532 54516 7534
rect 54908 9884 54964 9940
rect 55580 9938 55636 9940
rect 55580 9886 55582 9938
rect 55582 9886 55634 9938
rect 55634 9886 55636 9938
rect 55580 9884 55636 9886
rect 55244 7644 55300 7700
rect 55692 7698 55748 7700
rect 55692 7646 55694 7698
rect 55694 7646 55746 7698
rect 55746 7646 55748 7698
rect 55692 7644 55748 7646
rect 56252 7644 56308 7700
rect 55356 7532 55412 7588
rect 54012 6636 54068 6692
rect 55356 5404 55412 5460
rect 41916 5068 41972 5124
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 22428 3666 22484 3668
rect 22428 3614 22430 3666
rect 22430 3614 22482 3666
rect 22482 3614 22484 3666
rect 22428 3612 22484 3614
rect 43932 5122 43988 5124
rect 43932 5070 43934 5122
rect 43934 5070 43986 5122
rect 43986 5070 43988 5122
rect 43932 5068 43988 5070
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 43372 3500 43428 3556
rect 43708 3612 43764 3668
rect 45612 3666 45668 3668
rect 45612 3614 45614 3666
rect 45614 3614 45666 3666
rect 45666 3614 45668 3666
rect 45612 3612 45668 3614
rect 44940 3554 44996 3556
rect 44940 3502 44942 3554
rect 44942 3502 44994 3554
rect 44994 3502 44996 3554
rect 44940 3500 44996 3502
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 8306 52108 8316 52164
rect 8372 52108 8876 52164
rect 8932 52108 9100 52164
rect 9156 52108 9166 52164
rect 4162 51884 4172 51940
rect 4228 51884 8428 51940
rect 8484 51884 8494 51940
rect 8530 51772 8540 51828
rect 8596 51772 9324 51828
rect 9380 51772 9390 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 8978 51324 8988 51380
rect 9044 51324 9772 51380
rect 9828 51324 14140 51380
rect 14196 51324 14206 51380
rect 52434 51212 52444 51268
rect 52500 51212 55132 51268
rect 55188 51212 55198 51268
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 2034 50652 2044 50708
rect 2100 50652 5068 50708
rect 5124 50652 5134 50708
rect 4274 50540 4284 50596
rect 4340 50540 4956 50596
rect 5012 50540 6524 50596
rect 6580 50540 6590 50596
rect 10098 50540 10108 50596
rect 10164 50540 12012 50596
rect 12068 50540 13244 50596
rect 13300 50540 14364 50596
rect 14420 50540 14430 50596
rect 13906 50428 13916 50484
rect 13972 50428 15820 50484
rect 15876 50428 15886 50484
rect 16594 50428 16604 50484
rect 16660 50428 17052 50484
rect 17108 50428 17948 50484
rect 18004 50428 18508 50484
rect 18564 50428 19628 50484
rect 19684 50428 19694 50484
rect 24434 50428 24444 50484
rect 24500 50428 25900 50484
rect 25956 50428 26236 50484
rect 26292 50428 27692 50484
rect 27748 50428 27758 50484
rect 33954 50428 33964 50484
rect 34020 50428 36316 50484
rect 36372 50428 37436 50484
rect 37492 50428 39452 50484
rect 39508 50428 40012 50484
rect 40068 50428 40348 50484
rect 40404 50428 40414 50484
rect 53330 50428 53340 50484
rect 53396 50428 54236 50484
rect 54292 50428 54302 50484
rect 37650 50316 37660 50372
rect 37716 50316 39676 50372
rect 39732 50316 39742 50372
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 7298 49980 7308 50036
rect 7364 49980 9884 50036
rect 9940 49980 9950 50036
rect 10770 49980 10780 50036
rect 10836 49980 11676 50036
rect 11732 49980 11742 50036
rect 12450 49980 12460 50036
rect 12516 49980 13692 50036
rect 13748 49980 13758 50036
rect 46610 49980 46620 50036
rect 46676 49980 47628 50036
rect 47684 49980 47694 50036
rect 8754 49868 8764 49924
rect 8820 49868 9772 49924
rect 9828 49868 9838 49924
rect 19954 49868 19964 49924
rect 20020 49868 20972 49924
rect 21028 49868 21980 49924
rect 22036 49868 22046 49924
rect 24882 49868 24892 49924
rect 24948 49868 25788 49924
rect 25844 49868 25854 49924
rect 44034 49868 44044 49924
rect 44100 49868 47740 49924
rect 47796 49868 47806 49924
rect 11890 49756 11900 49812
rect 11956 49756 12684 49812
rect 12740 49756 12750 49812
rect 36866 49756 36876 49812
rect 36932 49756 42252 49812
rect 42308 49756 42318 49812
rect 42802 49756 42812 49812
rect 42868 49756 43932 49812
rect 43988 49756 43998 49812
rect 45938 49756 45948 49812
rect 46004 49756 46956 49812
rect 47012 49756 48972 49812
rect 49028 49756 49532 49812
rect 49588 49756 51100 49812
rect 51156 49756 53004 49812
rect 53060 49756 53564 49812
rect 53620 49756 53630 49812
rect 25106 49644 25116 49700
rect 25172 49644 25676 49700
rect 25732 49644 25742 49700
rect 26450 49644 26460 49700
rect 26516 49644 27356 49700
rect 27412 49644 27422 49700
rect 43250 49644 43260 49700
rect 43316 49644 44044 49700
rect 44100 49644 44110 49700
rect 10098 49532 10108 49588
rect 10164 49532 11564 49588
rect 11620 49532 13580 49588
rect 13636 49532 13646 49588
rect 24210 49532 24220 49588
rect 24276 49532 24780 49588
rect 24836 49532 26684 49588
rect 26740 49532 26750 49588
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 59200 49140 59800 49168
rect 20738 49084 20748 49140
rect 20804 49084 21868 49140
rect 21924 49084 21934 49140
rect 22978 49084 22988 49140
rect 23044 49084 24892 49140
rect 24948 49084 24958 49140
rect 55346 49084 55356 49140
rect 55412 49084 59800 49140
rect 59200 49056 59800 49084
rect 7298 48972 7308 49028
rect 7364 48972 8540 49028
rect 8596 48972 8606 49028
rect 17266 48972 17276 49028
rect 17332 48972 21644 49028
rect 21700 48972 21710 49028
rect 25106 48860 25116 48916
rect 25172 48860 26572 48916
rect 26628 48860 26638 48916
rect 28690 48860 28700 48916
rect 28756 48860 30044 48916
rect 30100 48860 30110 48916
rect 44706 48860 44716 48916
rect 44772 48860 45500 48916
rect 45556 48860 45566 48916
rect 48962 48860 48972 48916
rect 49028 48860 50316 48916
rect 50372 48860 50382 48916
rect 54338 48860 54348 48916
rect 54404 48860 56924 48916
rect 56980 48860 56990 48916
rect 7970 48748 7980 48804
rect 8036 48748 8652 48804
rect 8708 48748 8718 48804
rect 12898 48748 12908 48804
rect 12964 48748 13132 48804
rect 13188 48748 13804 48804
rect 13860 48748 14028 48804
rect 14084 48748 14094 48804
rect 33842 48748 33852 48804
rect 33908 48748 34412 48804
rect 34468 48748 34478 48804
rect 7522 48636 7532 48692
rect 7588 48636 8316 48692
rect 8372 48636 8764 48692
rect 8820 48636 8830 48692
rect 27010 48636 27020 48692
rect 27076 48636 27804 48692
rect 27860 48636 27870 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 24658 48412 24668 48468
rect 24724 48412 25564 48468
rect 25620 48412 26012 48468
rect 26068 48412 26078 48468
rect 4946 48300 4956 48356
rect 5012 48300 7308 48356
rect 7364 48300 7374 48356
rect 23202 48300 23212 48356
rect 23268 48300 24444 48356
rect 24500 48300 24510 48356
rect 7410 48188 7420 48244
rect 7476 48188 8988 48244
rect 9044 48188 9660 48244
rect 9716 48188 9726 48244
rect 12450 48188 12460 48244
rect 12516 48188 12796 48244
rect 12852 48188 13244 48244
rect 13300 48188 13916 48244
rect 13972 48188 13982 48244
rect 23426 48188 23436 48244
rect 23492 48188 24332 48244
rect 24388 48188 24398 48244
rect 48738 48188 48748 48244
rect 48804 48188 49532 48244
rect 49588 48188 50876 48244
rect 50932 48188 50942 48244
rect 10770 48076 10780 48132
rect 10836 48076 12908 48132
rect 12964 48076 12974 48132
rect 25666 48076 25676 48132
rect 25732 48076 26348 48132
rect 26404 48076 26414 48132
rect 40786 48076 40796 48132
rect 40852 48076 42476 48132
rect 42532 48076 42542 48132
rect 43026 48076 43036 48132
rect 43092 48076 43708 48132
rect 43764 48076 44492 48132
rect 44548 48076 44558 48132
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 21634 47628 21644 47684
rect 21700 47628 23212 47684
rect 23268 47628 23278 47684
rect 36530 47628 36540 47684
rect 36596 47628 37772 47684
rect 37828 47628 37838 47684
rect 7858 47516 7868 47572
rect 7924 47516 8652 47572
rect 8708 47516 8718 47572
rect 24322 47516 24332 47572
rect 24388 47516 25676 47572
rect 25732 47516 25742 47572
rect 36754 47516 36764 47572
rect 36820 47516 37996 47572
rect 38052 47516 38062 47572
rect 50082 47516 50092 47572
rect 50148 47516 53452 47572
rect 53508 47516 53518 47572
rect 28690 47404 28700 47460
rect 28756 47404 30268 47460
rect 30324 47404 30716 47460
rect 30772 47404 32172 47460
rect 32228 47404 32508 47460
rect 32564 47404 32574 47460
rect 52434 47404 52444 47460
rect 52500 47404 54012 47460
rect 54068 47404 54078 47460
rect 27794 47292 27804 47348
rect 27860 47292 28476 47348
rect 28532 47292 29484 47348
rect 29540 47292 29550 47348
rect 30930 47292 30940 47348
rect 30996 47292 31836 47348
rect 31892 47292 31902 47348
rect 44482 47292 44492 47348
rect 44548 47292 45612 47348
rect 45668 47292 45678 47348
rect 7634 47180 7644 47236
rect 7700 47180 8428 47236
rect 8484 47180 8764 47236
rect 8820 47180 10220 47236
rect 10276 47180 11900 47236
rect 11956 47180 11966 47236
rect 29810 47180 29820 47236
rect 29876 47180 31948 47236
rect 32004 47180 32014 47236
rect 45826 47180 45836 47236
rect 45892 47180 47180 47236
rect 47236 47180 47516 47236
rect 47572 47180 47582 47236
rect 7298 47068 7308 47124
rect 7364 47068 8316 47124
rect 8372 47068 8708 47124
rect 41570 47068 41580 47124
rect 41636 47068 42700 47124
rect 42756 47068 42766 47124
rect 52658 47068 52668 47124
rect 52724 47068 52734 47124
rect 8652 47012 8708 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 52668 47012 52724 47068
rect 8642 46956 8652 47012
rect 8708 46956 8718 47012
rect 38322 46956 38332 47012
rect 38388 46956 41692 47012
rect 41748 46956 41758 47012
rect 51538 46956 51548 47012
rect 51604 46956 54572 47012
rect 54628 46956 54638 47012
rect 16818 46844 16828 46900
rect 16884 46844 17612 46900
rect 17668 46844 17678 46900
rect 5730 46732 5740 46788
rect 5796 46732 8988 46788
rect 9044 46732 9054 46788
rect 14130 46732 14140 46788
rect 14196 46732 15036 46788
rect 15092 46732 16940 46788
rect 16996 46732 18396 46788
rect 18452 46732 18462 46788
rect 48402 46732 48412 46788
rect 48468 46732 54012 46788
rect 54068 46732 54078 46788
rect 9874 46620 9884 46676
rect 9940 46620 12012 46676
rect 12068 46620 12908 46676
rect 12964 46620 12974 46676
rect 26898 46620 26908 46676
rect 26964 46620 27468 46676
rect 27524 46620 27534 46676
rect 27682 46620 27692 46676
rect 27748 46620 28476 46676
rect 28532 46620 28542 46676
rect 42354 46620 42364 46676
rect 42420 46620 42700 46676
rect 42756 46620 42766 46676
rect 50418 46620 50428 46676
rect 50484 46620 51212 46676
rect 51268 46620 51548 46676
rect 51604 46620 51614 46676
rect 13682 46508 13692 46564
rect 13748 46508 15372 46564
rect 15428 46508 15438 46564
rect 24770 46508 24780 46564
rect 24836 46508 26124 46564
rect 26180 46508 26190 46564
rect 31266 46508 31276 46564
rect 31332 46508 32732 46564
rect 32788 46508 32798 46564
rect 47730 46508 47740 46564
rect 47796 46508 49532 46564
rect 49588 46508 54684 46564
rect 54740 46508 54750 46564
rect 42578 46396 42588 46452
rect 42644 46396 47068 46452
rect 47124 46396 47134 46452
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 17378 46060 17388 46116
rect 17444 46060 21756 46116
rect 21812 46060 21822 46116
rect 2818 45948 2828 46004
rect 2884 45948 3500 46004
rect 3556 45948 3566 46004
rect 4946 45948 4956 46004
rect 5012 45948 5404 46004
rect 5460 45948 5470 46004
rect 13570 45948 13580 46004
rect 13636 45948 14140 46004
rect 14196 45948 14206 46004
rect 20850 45948 20860 46004
rect 20916 45948 21868 46004
rect 21924 45948 21934 46004
rect 30818 45948 30828 46004
rect 30884 45948 31276 46004
rect 31332 45948 31342 46004
rect 46946 45948 46956 46004
rect 47012 45948 48972 46004
rect 49028 45948 50428 46004
rect 50484 45948 50494 46004
rect 12898 45836 12908 45892
rect 12964 45836 13916 45892
rect 13972 45836 14476 45892
rect 14532 45836 16828 45892
rect 16884 45836 17164 45892
rect 17220 45836 17230 45892
rect 24658 45836 24668 45892
rect 24724 45836 26796 45892
rect 26852 45836 27916 45892
rect 27972 45836 27982 45892
rect 37650 45836 37660 45892
rect 37716 45836 40796 45892
rect 40852 45836 41020 45892
rect 41076 45836 41468 45892
rect 41524 45836 43820 45892
rect 43876 45836 43886 45892
rect 5058 45612 5068 45668
rect 5124 45612 5628 45668
rect 5684 45612 5852 45668
rect 5908 45612 8092 45668
rect 8148 45612 8158 45668
rect 29810 45612 29820 45668
rect 29876 45612 32956 45668
rect 33012 45612 33022 45668
rect 42018 45612 42028 45668
rect 42084 45612 42364 45668
rect 42420 45612 42430 45668
rect 30594 45500 30604 45556
rect 30660 45500 31388 45556
rect 31444 45500 31454 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 16370 45388 16380 45444
rect 16436 45388 18060 45444
rect 18116 45388 18126 45444
rect 20178 45388 20188 45444
rect 20244 45388 21644 45444
rect 21700 45388 23212 45444
rect 23268 45388 23278 45444
rect 27906 45388 27916 45444
rect 27972 45388 28140 45444
rect 28196 45388 28476 45444
rect 28532 45388 31164 45444
rect 31220 45388 31724 45444
rect 31780 45388 31790 45444
rect 42018 45388 42028 45444
rect 42084 45388 43932 45444
rect 43988 45388 43998 45444
rect 15250 45276 15260 45332
rect 15316 45276 17724 45332
rect 17780 45276 17790 45332
rect 24098 45276 24108 45332
rect 24164 45276 26684 45332
rect 26740 45276 28812 45332
rect 28868 45276 28878 45332
rect 40786 45276 40796 45332
rect 40852 45276 41804 45332
rect 41860 45276 41870 45332
rect 25554 45164 25564 45220
rect 25620 45164 28196 45220
rect 28140 45108 28196 45164
rect 9874 45052 9884 45108
rect 9940 45052 10444 45108
rect 10500 45052 10510 45108
rect 25890 45052 25900 45108
rect 25956 45052 26236 45108
rect 26292 45052 26908 45108
rect 28130 45052 28140 45108
rect 28196 45052 30268 45108
rect 30324 45052 30334 45108
rect 40450 45052 40460 45108
rect 40516 45052 41580 45108
rect 41636 45052 41646 45108
rect 26852 44996 26908 45052
rect 26852 44940 28364 44996
rect 28420 44940 29708 44996
rect 29764 44940 29774 44996
rect 38098 44940 38108 44996
rect 38164 44940 41804 44996
rect 41860 44940 41870 44996
rect 46610 44940 46620 44996
rect 46676 44940 47404 44996
rect 47460 44940 47470 44996
rect 55122 44940 55132 44996
rect 55188 44940 55916 44996
rect 55972 44940 55982 44996
rect 24658 44828 24668 44884
rect 24724 44828 25788 44884
rect 25844 44828 26068 44884
rect 26012 44772 26068 44828
rect 26002 44716 26012 44772
rect 26068 44716 26078 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 25452 44604 26908 44660
rect 26964 44604 26974 44660
rect 25452 44548 25508 44604
rect 24882 44492 24892 44548
rect 24948 44492 25452 44548
rect 25508 44492 25518 44548
rect 26114 44492 26124 44548
rect 26180 44492 27244 44548
rect 27300 44492 27310 44548
rect 28914 44380 28924 44436
rect 28980 44380 29932 44436
rect 29988 44380 29998 44436
rect 5842 44268 5852 44324
rect 5908 44268 6412 44324
rect 6468 44268 6478 44324
rect 9986 44268 9996 44324
rect 10052 44268 10332 44324
rect 10388 44268 10398 44324
rect 20850 44268 20860 44324
rect 20916 44268 21756 44324
rect 21812 44268 21822 44324
rect 30146 44268 30156 44324
rect 30212 44268 30828 44324
rect 30884 44268 30894 44324
rect 52434 44268 52444 44324
rect 52500 44268 54012 44324
rect 54068 44268 54078 44324
rect 22530 44156 22540 44212
rect 22596 44156 26796 44212
rect 26852 44156 26862 44212
rect 48402 44156 48412 44212
rect 48468 44156 48972 44212
rect 49028 44156 49038 44212
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 200 43764 800 43792
rect 200 43708 4172 43764
rect 4228 43708 4238 43764
rect 48402 43708 48412 43764
rect 48468 43708 51100 43764
rect 51156 43708 51166 43764
rect 200 43680 800 43708
rect 52322 43596 52332 43652
rect 52388 43596 53004 43652
rect 53060 43596 53340 43652
rect 53396 43596 56252 43652
rect 56308 43596 56318 43652
rect 9314 43484 9324 43540
rect 9380 43484 10220 43540
rect 10276 43484 10286 43540
rect 18050 43484 18060 43540
rect 18116 43484 18396 43540
rect 18452 43484 18844 43540
rect 18900 43484 20188 43540
rect 20244 43484 20254 43540
rect 40226 43484 40236 43540
rect 40292 43484 42140 43540
rect 42196 43484 42476 43540
rect 42532 43484 42542 43540
rect 8306 43372 8316 43428
rect 8372 43372 10780 43428
rect 10836 43372 15036 43428
rect 15092 43372 15102 43428
rect 21186 43372 21196 43428
rect 21252 43372 22092 43428
rect 22148 43372 22158 43428
rect 49410 43372 49420 43428
rect 49476 43372 50876 43428
rect 50932 43372 51212 43428
rect 51268 43372 51278 43428
rect 6178 43260 6188 43316
rect 6244 43260 9884 43316
rect 9940 43260 9950 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 10098 42924 10108 42980
rect 10164 42924 14252 42980
rect 14308 42924 14318 42980
rect 14578 42924 14588 42980
rect 14644 42924 16044 42980
rect 16100 42924 16110 42980
rect 12898 42812 12908 42868
rect 12964 42812 15484 42868
rect 15540 42812 15550 42868
rect 23538 42812 23548 42868
rect 23604 42812 26124 42868
rect 26180 42812 26190 42868
rect 41570 42812 41580 42868
rect 41636 42812 42364 42868
rect 42420 42812 42430 42868
rect 14802 42700 14812 42756
rect 14868 42700 15596 42756
rect 15652 42700 15662 42756
rect 40674 42700 40684 42756
rect 40740 42700 42252 42756
rect 42308 42700 42318 42756
rect 43810 42700 43820 42756
rect 43876 42700 44716 42756
rect 44772 42700 44940 42756
rect 44996 42700 45612 42756
rect 45668 42700 46956 42756
rect 47012 42700 47022 42756
rect 50866 42700 50876 42756
rect 50932 42700 51884 42756
rect 51940 42700 51950 42756
rect 42802 42588 42812 42644
rect 42868 42588 44492 42644
rect 44548 42588 44558 42644
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 16482 42140 16492 42196
rect 16548 42140 17500 42196
rect 17556 42140 17566 42196
rect 25778 42140 25788 42196
rect 25844 42140 26572 42196
rect 26628 42140 27804 42196
rect 27860 42140 27870 42196
rect 53330 42140 53340 42196
rect 53396 42140 54124 42196
rect 54180 42140 54190 42196
rect 31602 42028 31612 42084
rect 31668 42028 33628 42084
rect 33684 42028 34748 42084
rect 34804 42028 35756 42084
rect 35812 42028 36988 42084
rect 37044 42028 38108 42084
rect 38164 42028 38174 42084
rect 39330 42028 39340 42084
rect 39396 42028 42588 42084
rect 42644 42028 42654 42084
rect 49634 42028 49644 42084
rect 49700 42028 50092 42084
rect 50148 42028 50876 42084
rect 50932 42028 50942 42084
rect 2146 41916 2156 41972
rect 2212 41916 4396 41972
rect 4452 41916 5852 41972
rect 5908 41916 5918 41972
rect 6066 41916 6076 41972
rect 6132 41916 8428 41972
rect 8484 41916 9324 41972
rect 9380 41916 9996 41972
rect 10052 41916 10332 41972
rect 10388 41916 11676 41972
rect 11732 41916 13580 41972
rect 13636 41916 13646 41972
rect 15026 41916 15036 41972
rect 15092 41916 15820 41972
rect 15876 41916 15886 41972
rect 19394 41916 19404 41972
rect 19460 41916 20300 41972
rect 20356 41916 20860 41972
rect 20916 41916 20926 41972
rect 26450 41916 26460 41972
rect 26516 41916 29260 41972
rect 29316 41916 29326 41972
rect 36530 41916 36540 41972
rect 36596 41916 38780 41972
rect 38836 41916 38846 41972
rect 5058 41804 5068 41860
rect 5124 41804 5628 41860
rect 5684 41804 5694 41860
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 32050 41356 32060 41412
rect 32116 41356 35196 41412
rect 35252 41356 35262 41412
rect 20626 41244 20636 41300
rect 20692 41244 21868 41300
rect 21924 41244 21934 41300
rect 34402 41244 34412 41300
rect 34468 41244 35308 41300
rect 35364 41244 35374 41300
rect 11666 41132 11676 41188
rect 11732 41132 12348 41188
rect 12404 41132 12414 41188
rect 17154 41132 17164 41188
rect 17220 41132 17724 41188
rect 17780 41132 19404 41188
rect 19460 41132 19470 41188
rect 10770 41020 10780 41076
rect 10836 41020 11788 41076
rect 11844 41020 11854 41076
rect 23202 41020 23212 41076
rect 23268 41020 26908 41076
rect 26964 41020 26974 41076
rect 42466 40908 42476 40964
rect 42532 40908 44380 40964
rect 44436 40908 46844 40964
rect 46900 40908 46910 40964
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 13010 40460 13020 40516
rect 13076 40460 13692 40516
rect 13748 40460 13758 40516
rect 19954 40460 19964 40516
rect 20020 40460 21644 40516
rect 21700 40460 21710 40516
rect 22978 40460 22988 40516
rect 23044 40460 24332 40516
rect 24388 40460 24398 40516
rect 28578 40460 28588 40516
rect 28644 40460 29260 40516
rect 29316 40460 29326 40516
rect 15026 40348 15036 40404
rect 15092 40348 19068 40404
rect 19124 40348 21084 40404
rect 21140 40348 26684 40404
rect 26740 40348 27244 40404
rect 27300 40348 27310 40404
rect 37874 40348 37884 40404
rect 37940 40348 38780 40404
rect 38836 40348 40908 40404
rect 40964 40348 40974 40404
rect 35634 40236 35644 40292
rect 35700 40236 37324 40292
rect 37380 40236 37390 40292
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 25666 39676 25676 39732
rect 25732 39676 27020 39732
rect 27076 39676 27086 39732
rect 46610 39676 46620 39732
rect 46676 39676 47628 39732
rect 47684 39676 49868 39732
rect 49924 39676 49934 39732
rect 53666 39676 53676 39732
rect 53732 39676 54572 39732
rect 54628 39676 54638 39732
rect 22306 39564 22316 39620
rect 22372 39564 24556 39620
rect 24612 39564 25564 39620
rect 25620 39564 27692 39620
rect 27748 39564 27758 39620
rect 29698 39564 29708 39620
rect 29764 39564 32172 39620
rect 32228 39564 32956 39620
rect 33012 39564 33022 39620
rect 46834 39564 46844 39620
rect 46900 39564 51212 39620
rect 51268 39564 52332 39620
rect 52388 39564 52398 39620
rect 47618 39452 47628 39508
rect 47684 39452 49532 39508
rect 49588 39452 53676 39508
rect 53732 39452 53742 39508
rect 20290 39340 20300 39396
rect 20356 39340 21532 39396
rect 21588 39340 22764 39396
rect 22820 39340 23548 39396
rect 23604 39340 23614 39396
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 49746 39116 49756 39172
rect 49812 39116 50092 39172
rect 50148 39116 50158 39172
rect 50092 39060 50148 39116
rect 43362 39004 43372 39060
rect 43428 39004 44044 39060
rect 44100 39004 44110 39060
rect 50092 39004 51212 39060
rect 51268 39004 51278 39060
rect 32834 38892 32844 38948
rect 32900 38892 33628 38948
rect 33684 38892 33694 38948
rect 52322 38892 52332 38948
rect 52388 38892 53452 38948
rect 53508 38892 53518 38948
rect 7746 38780 7756 38836
rect 7812 38780 9772 38836
rect 9828 38780 9838 38836
rect 25106 38780 25116 38836
rect 25172 38780 26796 38836
rect 26852 38780 26862 38836
rect 27682 38780 27692 38836
rect 27748 38780 28364 38836
rect 28420 38780 31612 38836
rect 31668 38780 31678 38836
rect 35074 38780 35084 38836
rect 35140 38780 40012 38836
rect 40068 38780 40078 38836
rect 43474 38780 43484 38836
rect 43540 38780 47572 38836
rect 47730 38780 47740 38836
rect 47796 38780 49532 38836
rect 49588 38780 49598 38836
rect 51650 38780 51660 38836
rect 51716 38780 52444 38836
rect 52500 38780 54012 38836
rect 54068 38780 54078 38836
rect 47516 38724 47572 38780
rect 36978 38668 36988 38724
rect 37044 38668 40348 38724
rect 40404 38668 40414 38724
rect 42802 38668 42812 38724
rect 42868 38668 44380 38724
rect 44436 38668 44446 38724
rect 47516 38668 48188 38724
rect 48244 38668 48254 38724
rect 50978 38668 50988 38724
rect 51044 38668 51436 38724
rect 51492 38668 53004 38724
rect 53060 38668 53070 38724
rect 53330 38668 53340 38724
rect 53396 38668 54124 38724
rect 54180 38668 54190 38724
rect 37650 38556 37660 38612
rect 37716 38556 39676 38612
rect 39732 38556 39742 38612
rect 48738 38556 48748 38612
rect 48804 38556 49756 38612
rect 49812 38556 49822 38612
rect 52882 38556 52892 38612
rect 52948 38556 54236 38612
rect 54292 38556 54302 38612
rect 48178 38444 48188 38500
rect 48244 38444 49980 38500
rect 50036 38444 50652 38500
rect 50708 38444 50718 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 12674 38108 12684 38164
rect 12740 38108 13356 38164
rect 13412 38108 15036 38164
rect 15092 38108 15102 38164
rect 34962 38108 34972 38164
rect 35028 38108 36316 38164
rect 36372 38108 36382 38164
rect 36642 38108 36652 38164
rect 36708 38108 37548 38164
rect 37604 38108 37614 38164
rect 52098 38108 52108 38164
rect 52164 38108 52780 38164
rect 52836 38108 54348 38164
rect 54404 38108 56364 38164
rect 56420 38108 56430 38164
rect 12684 38052 12740 38108
rect 8306 37996 8316 38052
rect 8372 37996 12740 38052
rect 14690 37996 14700 38052
rect 14756 37996 15484 38052
rect 15540 37996 15550 38052
rect 36754 37884 36764 37940
rect 36820 37884 37884 37940
rect 37940 37884 37950 37940
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 7858 37436 7868 37492
rect 7924 37436 8764 37492
rect 8820 37436 10892 37492
rect 10948 37436 11228 37492
rect 11284 37436 11788 37492
rect 11844 37436 11854 37492
rect 24210 37436 24220 37492
rect 24276 37436 26684 37492
rect 26740 37436 26750 37492
rect 38322 37436 38332 37492
rect 38388 37436 42924 37492
rect 42980 37436 42990 37492
rect 34626 37324 34636 37380
rect 34692 37324 35532 37380
rect 35588 37324 35598 37380
rect 52546 37324 52556 37380
rect 52612 37324 53676 37380
rect 53732 37324 53742 37380
rect 32162 37212 32172 37268
rect 32228 37212 33852 37268
rect 33908 37212 35084 37268
rect 35140 37212 36988 37268
rect 37044 37212 37054 37268
rect 48402 37212 48412 37268
rect 48468 37212 48972 37268
rect 49028 37212 49532 37268
rect 49588 37212 49598 37268
rect 49746 37212 49756 37268
rect 49812 37212 51324 37268
rect 51380 37212 51390 37268
rect 51538 37212 51548 37268
rect 51604 37212 53564 37268
rect 53620 37212 53630 37268
rect 51324 37156 51380 37212
rect 32498 37100 32508 37156
rect 32564 37100 37436 37156
rect 37492 37100 37502 37156
rect 47842 37100 47852 37156
rect 47908 37100 48468 37156
rect 51324 37100 52108 37156
rect 52164 37100 52174 37156
rect 48412 37044 48468 37100
rect 31490 36988 31500 37044
rect 31556 36988 32172 37044
rect 32228 36988 32238 37044
rect 46946 36988 46956 37044
rect 47012 36988 48076 37044
rect 48132 36988 48142 37044
rect 48402 36988 48412 37044
rect 48468 36988 50092 37044
rect 50148 36988 50158 37044
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 7746 36652 7756 36708
rect 7812 36652 8316 36708
rect 8372 36652 8382 36708
rect 7970 36540 7980 36596
rect 8036 36540 9100 36596
rect 9156 36540 9166 36596
rect 16146 36540 16156 36596
rect 16212 36540 17388 36596
rect 17444 36540 17454 36596
rect 24882 36540 24892 36596
rect 24948 36540 25340 36596
rect 25396 36540 25406 36596
rect 36978 36540 36988 36596
rect 37044 36540 37548 36596
rect 37604 36540 37614 36596
rect 43474 36540 43484 36596
rect 43540 36540 46284 36596
rect 46340 36540 46844 36596
rect 46900 36540 46910 36596
rect 40786 36428 40796 36484
rect 40852 36428 43148 36484
rect 43204 36428 43214 36484
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 4498 35644 4508 35700
rect 4564 35644 5404 35700
rect 5460 35644 7756 35700
rect 7812 35644 7822 35700
rect 12450 35644 12460 35700
rect 12516 35644 13244 35700
rect 13300 35644 14476 35700
rect 14532 35644 16604 35700
rect 16660 35644 17612 35700
rect 17668 35644 17948 35700
rect 18004 35644 18284 35700
rect 18340 35644 18350 35700
rect 21186 35644 21196 35700
rect 21252 35644 23548 35700
rect 23604 35644 24444 35700
rect 24500 35644 24510 35700
rect 27906 35644 27916 35700
rect 27972 35644 28588 35700
rect 28644 35644 31948 35700
rect 32004 35644 32014 35700
rect 22978 35532 22988 35588
rect 23044 35532 23996 35588
rect 24052 35532 24062 35588
rect 33058 35532 33068 35588
rect 33124 35532 36092 35588
rect 36148 35532 36158 35588
rect 41794 35308 41804 35364
rect 41860 35308 43596 35364
rect 43652 35308 43662 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 39442 35196 39452 35252
rect 39508 35196 40572 35252
rect 40628 35196 41468 35252
rect 41524 35196 44716 35252
rect 44772 35196 44782 35252
rect 20850 35084 20860 35140
rect 20916 35084 22428 35140
rect 22484 35084 22494 35140
rect 13682 34860 13692 34916
rect 13748 34860 14252 34916
rect 14308 34860 15036 34916
rect 15092 34860 15102 34916
rect 44706 34860 44716 34916
rect 44772 34860 45276 34916
rect 45332 34860 45342 34916
rect 8194 34748 8204 34804
rect 8260 34748 8988 34804
rect 9044 34748 9054 34804
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 46834 34300 46844 34356
rect 46900 34300 47740 34356
rect 47796 34300 47806 34356
rect 16482 34188 16492 34244
rect 16548 34188 17724 34244
rect 17780 34188 17790 34244
rect 36530 34188 36540 34244
rect 36596 34188 37436 34244
rect 37492 34188 37502 34244
rect 15474 34076 15484 34132
rect 15540 34076 16716 34132
rect 16772 34076 18732 34132
rect 18788 34076 18798 34132
rect 38210 34076 38220 34132
rect 38276 34076 39452 34132
rect 39508 34076 39518 34132
rect 41346 34076 41356 34132
rect 41412 34076 41916 34132
rect 41972 34076 41982 34132
rect 6178 33964 6188 34020
rect 6244 33964 9772 34020
rect 9828 33964 12236 34020
rect 12292 33964 12302 34020
rect 35298 33964 35308 34020
rect 35364 33964 36428 34020
rect 36484 33964 36494 34020
rect 45378 33964 45388 34020
rect 45444 33964 46284 34020
rect 46340 33964 48076 34020
rect 48132 33964 48142 34020
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 20738 33628 20748 33684
rect 20804 33628 22428 33684
rect 22484 33628 22494 33684
rect 40562 33628 40572 33684
rect 40628 33628 41580 33684
rect 41636 33628 42812 33684
rect 42868 33628 42878 33684
rect 36530 33292 36540 33348
rect 36596 33292 37660 33348
rect 37716 33292 37726 33348
rect 36306 33068 36316 33124
rect 36372 33068 36764 33124
rect 36820 33068 37660 33124
rect 37716 33068 37726 33124
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 12898 32732 12908 32788
rect 12964 32732 13804 32788
rect 13860 32732 16156 32788
rect 16212 32732 17164 32788
rect 17220 32732 17230 32788
rect 32722 32620 32732 32676
rect 32788 32620 33628 32676
rect 33684 32620 33694 32676
rect 24882 32396 24892 32452
rect 24948 32396 27020 32452
rect 27076 32396 27086 32452
rect 43810 32396 43820 32452
rect 43876 32396 44940 32452
rect 44996 32396 45612 32452
rect 45668 32396 46172 32452
rect 46228 32396 46238 32452
rect 34738 32284 34748 32340
rect 34804 32284 35980 32340
rect 36036 32284 36046 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 14354 31836 14364 31892
rect 14420 31836 15708 31892
rect 15764 31836 15774 31892
rect 17938 31836 17948 31892
rect 18004 31836 19404 31892
rect 19460 31836 19628 31892
rect 19684 31836 20860 31892
rect 20916 31836 20926 31892
rect 45378 31724 45388 31780
rect 45444 31724 46844 31780
rect 46900 31724 51212 31780
rect 51268 31724 51278 31780
rect 19282 31500 19292 31556
rect 19348 31500 20300 31556
rect 20356 31500 20366 31556
rect 31938 31500 31948 31556
rect 32004 31500 32508 31556
rect 32564 31500 33740 31556
rect 33796 31500 35196 31556
rect 35252 31500 35262 31556
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 12898 31164 12908 31220
rect 12964 31164 16268 31220
rect 16324 31164 16334 31220
rect 5954 31052 5964 31108
rect 6020 31052 6188 31108
rect 6244 31052 6412 31108
rect 6468 31052 10108 31108
rect 10164 31052 10174 31108
rect 36754 31052 36764 31108
rect 36820 31052 37884 31108
rect 37940 31052 37950 31108
rect 15026 30940 15036 30996
rect 15092 30940 15372 30996
rect 15428 30940 18508 30996
rect 18564 30940 19068 30996
rect 19124 30940 19134 30996
rect 29698 30940 29708 30996
rect 29764 30940 29932 30996
rect 29988 30940 31948 30996
rect 32004 30940 32014 30996
rect 45938 30940 45948 30996
rect 46004 30940 49532 30996
rect 49588 30940 49598 30996
rect 3042 30828 3052 30884
rect 3108 30828 5068 30884
rect 5124 30828 5134 30884
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19170 30380 19180 30436
rect 19236 30380 20188 30436
rect 20244 30380 20254 30436
rect 49746 30380 49756 30436
rect 49812 30380 52444 30436
rect 52500 30380 52510 30436
rect 16370 30268 16380 30324
rect 16436 30268 16716 30324
rect 16772 30268 18620 30324
rect 18676 30268 20300 30324
rect 20356 30268 21644 30324
rect 21700 30268 21710 30324
rect 32274 30268 32284 30324
rect 32340 30268 32732 30324
rect 32788 30268 33292 30324
rect 33348 30268 33358 30324
rect 39666 30268 39676 30324
rect 39732 30268 40236 30324
rect 40292 30268 40302 30324
rect 48514 30268 48524 30324
rect 48580 30268 49532 30324
rect 49588 30268 49598 30324
rect 20066 30156 20076 30212
rect 20132 30156 20524 30212
rect 20580 30156 20590 30212
rect 37650 30156 37660 30212
rect 37716 30156 38556 30212
rect 38612 30156 44156 30212
rect 44212 30156 45388 30212
rect 45444 30156 45454 30212
rect 36978 30044 36988 30100
rect 37044 30044 40348 30100
rect 40404 30044 40796 30100
rect 40852 30044 40862 30100
rect 27234 29932 27244 29988
rect 27300 29932 28140 29988
rect 28196 29932 28206 29988
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 12226 29596 12236 29652
rect 12292 29596 13132 29652
rect 13188 29596 13198 29652
rect 8978 29372 8988 29428
rect 9044 29372 9660 29428
rect 9716 29372 9726 29428
rect 24098 29372 24108 29428
rect 24164 29372 26572 29428
rect 26628 29372 27356 29428
rect 27412 29372 28140 29428
rect 28196 29372 28206 29428
rect 33730 29372 33740 29428
rect 33796 29372 36988 29428
rect 37044 29372 37054 29428
rect 40786 29372 40796 29428
rect 40852 29372 41580 29428
rect 41636 29372 41646 29428
rect 36530 29260 36540 29316
rect 36596 29260 39116 29316
rect 39172 29260 39182 29316
rect 44482 29260 44492 29316
rect 44548 29260 45388 29316
rect 45444 29260 45454 29316
rect 45938 29260 45948 29316
rect 46004 29260 49532 29316
rect 49588 29260 49598 29316
rect 38210 29148 38220 29204
rect 38276 29148 39228 29204
rect 39284 29148 39294 29204
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 6626 28812 6636 28868
rect 6692 28812 7532 28868
rect 7588 28812 8204 28868
rect 8260 28812 8270 28868
rect 24882 28812 24892 28868
rect 24948 28812 25900 28868
rect 25956 28812 25966 28868
rect 4162 28700 4172 28756
rect 4228 28700 8428 28756
rect 18722 28700 18732 28756
rect 18788 28700 33404 28756
rect 33460 28700 34972 28756
rect 35028 28700 41356 28756
rect 41412 28700 41422 28756
rect 8372 28644 8428 28700
rect 5170 28588 5180 28644
rect 5236 28588 6188 28644
rect 6244 28588 6254 28644
rect 8372 28588 28252 28644
rect 28308 28588 30268 28644
rect 30324 28588 30334 28644
rect 5394 28476 5404 28532
rect 5460 28476 5964 28532
rect 6020 28476 7308 28532
rect 7364 28476 7374 28532
rect 19506 28476 19516 28532
rect 19572 28476 20412 28532
rect 20468 28476 20478 28532
rect 9426 28364 9436 28420
rect 9492 28364 15148 28420
rect 15204 28364 15214 28420
rect 21186 28364 21196 28420
rect 21252 28364 25788 28420
rect 25844 28364 25854 28420
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 15698 28028 15708 28084
rect 15764 28028 21756 28084
rect 21812 28028 21822 28084
rect 26338 28028 26348 28084
rect 26404 28028 27692 28084
rect 27748 28028 27758 28084
rect 21522 27916 21532 27972
rect 21588 27916 26236 27972
rect 26292 27916 26302 27972
rect 24994 27804 25004 27860
rect 25060 27804 25676 27860
rect 25732 27804 26348 27860
rect 26404 27804 26414 27860
rect 29362 27804 29372 27860
rect 29428 27804 31500 27860
rect 31556 27804 31566 27860
rect 43474 27804 43484 27860
rect 43540 27804 46508 27860
rect 46564 27804 46732 27860
rect 46788 27804 48076 27860
rect 48132 27804 49756 27860
rect 49812 27804 52108 27860
rect 52164 27804 53340 27860
rect 53396 27804 53406 27860
rect 14914 27692 14924 27748
rect 14980 27692 16380 27748
rect 16436 27692 16446 27748
rect 31378 27580 31388 27636
rect 31444 27580 31948 27636
rect 32004 27580 32014 27636
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 12898 27356 12908 27412
rect 12964 27356 14700 27412
rect 14756 27356 14766 27412
rect 15026 27244 15036 27300
rect 15092 27244 15820 27300
rect 15876 27244 15886 27300
rect 12898 27132 12908 27188
rect 12964 27132 14812 27188
rect 14868 27132 14878 27188
rect 35074 27020 35084 27076
rect 35140 27020 35756 27076
rect 35812 27020 37884 27076
rect 37940 27020 37950 27076
rect 39778 27020 39788 27076
rect 39844 27020 41804 27076
rect 41860 27020 41870 27076
rect 50204 27020 51660 27076
rect 51716 27020 51726 27076
rect 10098 26908 10108 26964
rect 10164 26908 11228 26964
rect 11284 26908 13020 26964
rect 13076 26908 13580 26964
rect 13636 26908 14924 26964
rect 14980 26908 14990 26964
rect 32274 26908 32284 26964
rect 32340 26908 34244 26964
rect 48514 26908 48524 26964
rect 48580 26908 49756 26964
rect 49812 26908 49822 26964
rect 6514 26796 6524 26852
rect 6580 26796 6860 26852
rect 6916 26796 7532 26852
rect 7588 26796 7598 26852
rect 34188 26740 34244 26908
rect 50204 26740 50260 27020
rect 59200 26964 59800 26992
rect 51538 26908 51548 26964
rect 51604 26908 52332 26964
rect 52388 26908 52398 26964
rect 55346 26908 55356 26964
rect 55412 26908 59800 26964
rect 59200 26880 59800 26908
rect 50642 26796 50652 26852
rect 50708 26796 53676 26852
rect 53732 26796 53742 26852
rect 34178 26684 34188 26740
rect 34244 26684 34254 26740
rect 50194 26684 50204 26740
rect 50260 26684 50270 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 23986 26460 23996 26516
rect 24052 26460 24892 26516
rect 24948 26460 25564 26516
rect 25620 26460 28140 26516
rect 28196 26460 28588 26516
rect 28644 26460 30492 26516
rect 30548 26460 31836 26516
rect 31892 26460 31902 26516
rect 42354 26460 42364 26516
rect 42420 26460 43708 26516
rect 7298 26348 7308 26404
rect 7364 26348 7980 26404
rect 8036 26348 9996 26404
rect 10052 26348 10062 26404
rect 40226 26236 40236 26292
rect 40292 26236 42812 26292
rect 42868 26236 42878 26292
rect 43652 26180 43708 26460
rect 47516 26348 48860 26404
rect 48916 26348 49644 26404
rect 49700 26348 49868 26404
rect 49924 26348 49934 26404
rect 50978 26348 50988 26404
rect 51044 26348 51324 26404
rect 51380 26348 51390 26404
rect 47516 26180 47572 26348
rect 48738 26236 48748 26292
rect 48804 26236 49532 26292
rect 49588 26236 49598 26292
rect 51090 26236 51100 26292
rect 51156 26236 51436 26292
rect 51492 26236 51502 26292
rect 4162 26124 4172 26180
rect 4228 26124 6188 26180
rect 6244 26124 6254 26180
rect 7522 26124 7532 26180
rect 7588 26124 9828 26180
rect 24434 26124 24444 26180
rect 24500 26124 26124 26180
rect 26180 26124 26190 26180
rect 40786 26124 40796 26180
rect 40852 26124 42028 26180
rect 42084 26124 42094 26180
rect 43652 26124 47516 26180
rect 47572 26124 47582 26180
rect 9772 26068 9828 26124
rect 7858 26012 7868 26068
rect 7924 26012 8764 26068
rect 8820 26012 8830 26068
rect 9762 26012 9772 26068
rect 9828 26012 9838 26068
rect 39778 26012 39788 26068
rect 39844 26012 41804 26068
rect 41860 26012 41870 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 6290 25676 6300 25732
rect 6356 25676 6972 25732
rect 7028 25676 8204 25732
rect 8260 25676 8270 25732
rect 18610 25564 18620 25620
rect 18676 25564 20300 25620
rect 20356 25564 20366 25620
rect 25106 25564 25116 25620
rect 25172 25564 25788 25620
rect 25844 25564 25854 25620
rect 49634 25564 49644 25620
rect 49700 25564 50428 25620
rect 50484 25564 50494 25620
rect 15810 25452 15820 25508
rect 15876 25452 17836 25508
rect 17892 25452 18284 25508
rect 18340 25452 18350 25508
rect 20178 25452 20188 25508
rect 20244 25452 20860 25508
rect 20916 25452 20926 25508
rect 21634 25452 21644 25508
rect 21700 25452 22316 25508
rect 22372 25452 23996 25508
rect 24052 25452 24062 25508
rect 31378 25452 31388 25508
rect 31444 25452 34748 25508
rect 34804 25452 34814 25508
rect 40114 25452 40124 25508
rect 40180 25452 41804 25508
rect 41860 25452 41870 25508
rect 48738 25452 48748 25508
rect 48804 25452 49868 25508
rect 49924 25452 49934 25508
rect 44706 25340 44716 25396
rect 44772 25340 45500 25396
rect 45556 25340 45566 25396
rect 49522 25340 49532 25396
rect 49588 25340 50876 25396
rect 50932 25340 50942 25396
rect 44482 25228 44492 25284
rect 44548 25228 45388 25284
rect 45444 25228 48076 25284
rect 48132 25228 48412 25284
rect 48468 25228 48478 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 16482 24892 16492 24948
rect 16548 24892 17724 24948
rect 17780 24892 17790 24948
rect 43652 24836 43708 24948
rect 43764 24892 44940 24948
rect 44996 24892 46844 24948
rect 46900 24892 46910 24948
rect 41794 24780 41804 24836
rect 41860 24780 43708 24836
rect 51202 24668 51212 24724
rect 51268 24668 51548 24724
rect 51604 24668 52444 24724
rect 52500 24668 52510 24724
rect 20738 24556 20748 24612
rect 20804 24556 21756 24612
rect 21812 24556 21822 24612
rect 42578 24556 42588 24612
rect 42644 24556 45612 24612
rect 45668 24556 45678 24612
rect 55346 24556 55356 24612
rect 55412 24556 55916 24612
rect 55972 24556 55982 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 52658 24108 52668 24164
rect 52724 24108 54572 24164
rect 54628 24108 54638 24164
rect 13010 23996 13020 24052
rect 13076 23996 17052 24052
rect 17108 23996 17118 24052
rect 24658 23996 24668 24052
rect 24724 23996 25676 24052
rect 25732 23996 25742 24052
rect 26786 23996 26796 24052
rect 26852 23996 29708 24052
rect 29764 23996 29774 24052
rect 44706 23996 44716 24052
rect 44772 23996 47068 24052
rect 47124 23996 47134 24052
rect 32162 23884 32172 23940
rect 32228 23884 34300 23940
rect 34356 23884 34366 23940
rect 36194 23884 36204 23940
rect 36260 23884 36540 23940
rect 36596 23884 37548 23940
rect 37604 23884 37614 23940
rect 12898 23772 12908 23828
rect 12964 23772 14476 23828
rect 14532 23772 14542 23828
rect 30370 23772 30380 23828
rect 30436 23772 31500 23828
rect 31556 23772 31566 23828
rect 17938 23660 17948 23716
rect 18004 23660 18284 23716
rect 18340 23660 18844 23716
rect 18900 23660 20188 23716
rect 20244 23660 20972 23716
rect 21028 23660 22204 23716
rect 22260 23660 22270 23716
rect 26674 23660 26684 23716
rect 26740 23660 27356 23716
rect 27412 23660 27422 23716
rect 31826 23660 31836 23716
rect 31892 23660 32844 23716
rect 32900 23660 32910 23716
rect 38658 23660 38668 23716
rect 38724 23660 41020 23716
rect 41076 23660 41086 23716
rect 47954 23660 47964 23716
rect 48020 23660 49532 23716
rect 49588 23660 51660 23716
rect 51716 23660 52556 23716
rect 52612 23660 52622 23716
rect 3948 23548 7084 23604
rect 7140 23548 7150 23604
rect 16594 23548 16604 23604
rect 16660 23548 18508 23604
rect 18564 23548 18574 23604
rect 32386 23548 32396 23604
rect 32452 23548 36764 23604
rect 36820 23548 36830 23604
rect 46386 23548 46396 23604
rect 46452 23548 46462 23604
rect 3948 23492 4004 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 46396 23492 46452 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 2706 23436 2716 23492
rect 2772 23436 3388 23492
rect 3444 23436 3454 23492
rect 3938 23436 3948 23492
rect 4004 23436 4014 23492
rect 46396 23436 47740 23492
rect 47796 23436 47806 23492
rect 46620 23380 46676 23436
rect 11218 23324 11228 23380
rect 11284 23324 11788 23380
rect 11844 23324 13020 23380
rect 13076 23324 13086 23380
rect 14578 23324 14588 23380
rect 14644 23324 14924 23380
rect 14980 23324 16604 23380
rect 16660 23324 16670 23380
rect 46610 23324 46620 23380
rect 46676 23324 46686 23380
rect 48066 23324 48076 23380
rect 48132 23324 51100 23380
rect 51156 23324 52220 23380
rect 52276 23324 52286 23380
rect 6066 23212 6076 23268
rect 6132 23212 6860 23268
rect 6916 23212 8428 23268
rect 8484 23212 9660 23268
rect 9716 23212 9726 23268
rect 13346 23212 13356 23268
rect 13412 23212 13804 23268
rect 13860 23212 13870 23268
rect 23426 23212 23436 23268
rect 23492 23212 26348 23268
rect 26404 23212 26908 23268
rect 12002 23100 12012 23156
rect 12068 23100 12684 23156
rect 12740 23100 13132 23156
rect 13188 23100 13580 23156
rect 13636 23100 13646 23156
rect 26852 23100 26908 23212
rect 26964 23100 26974 23156
rect 42018 23100 42028 23156
rect 42084 23100 42812 23156
rect 42868 23100 42878 23156
rect 48290 23100 48300 23156
rect 48356 23100 49756 23156
rect 49812 23100 50988 23156
rect 51044 23100 51054 23156
rect 51762 23100 51772 23156
rect 51828 23100 52780 23156
rect 52836 23100 52846 23156
rect 6626 22988 6636 23044
rect 6692 22988 11228 23044
rect 11284 22988 11294 23044
rect 27682 22988 27692 23044
rect 27748 22988 28924 23044
rect 28980 22988 28990 23044
rect 33618 22988 33628 23044
rect 33684 22988 34860 23044
rect 34916 22988 34926 23044
rect 50418 22876 50428 22932
rect 50484 22876 51548 22932
rect 51604 22876 52556 22932
rect 52612 22876 52622 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 33954 22652 33964 22708
rect 34020 22652 34972 22708
rect 35028 22652 35038 22708
rect 47394 22652 47404 22708
rect 47460 22652 48076 22708
rect 48132 22652 48142 22708
rect 47170 22540 47180 22596
rect 47236 22540 48300 22596
rect 48356 22540 48366 22596
rect 8418 22428 8428 22484
rect 8484 22428 8988 22484
rect 9044 22428 9054 22484
rect 15250 22428 15260 22484
rect 15316 22428 16044 22484
rect 16100 22428 16110 22484
rect 17378 22428 17388 22484
rect 17444 22428 18060 22484
rect 18116 22428 18126 22484
rect 9090 22316 9100 22372
rect 9156 22316 12012 22372
rect 12068 22316 12078 22372
rect 26002 22316 26012 22372
rect 26068 22316 27692 22372
rect 27748 22316 27758 22372
rect 37986 22316 37996 22372
rect 38052 22316 39228 22372
rect 39284 22316 39294 22372
rect 45602 22316 45612 22372
rect 45668 22316 46284 22372
rect 46340 22316 46350 22372
rect 47058 22316 47068 22372
rect 47124 22316 47964 22372
rect 48020 22316 48030 22372
rect 51090 22316 51100 22372
rect 51156 22316 51436 22372
rect 51492 22316 51502 22372
rect 34626 22204 34636 22260
rect 34692 22204 35756 22260
rect 35812 22204 35822 22260
rect 45826 22204 45836 22260
rect 45892 22204 46508 22260
rect 46564 22204 46574 22260
rect 46060 21980 48076 22036
rect 48132 21980 48142 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 46060 21924 46116 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 2258 21868 2268 21924
rect 2324 21868 2716 21924
rect 2772 21868 4732 21924
rect 4788 21868 4956 21924
rect 5012 21868 5628 21924
rect 5684 21868 6076 21924
rect 6132 21868 6142 21924
rect 46050 21868 46060 21924
rect 46116 21868 46126 21924
rect 47170 21868 47180 21924
rect 47236 21868 49644 21924
rect 49700 21868 50372 21924
rect 50316 21812 50372 21868
rect 50316 21756 50876 21812
rect 50932 21756 51436 21812
rect 51492 21756 51502 21812
rect 23202 21644 23212 21700
rect 23268 21644 25676 21700
rect 25732 21644 25742 21700
rect 32946 21644 32956 21700
rect 33012 21644 33740 21700
rect 33796 21644 35084 21700
rect 35140 21644 35644 21700
rect 35700 21644 35710 21700
rect 39218 21644 39228 21700
rect 39284 21644 41468 21700
rect 41524 21644 42140 21700
rect 42196 21644 42206 21700
rect 200 21588 800 21616
rect 200 21532 2492 21588
rect 2548 21532 2558 21588
rect 9426 21532 9436 21588
rect 9492 21532 9884 21588
rect 9940 21532 13132 21588
rect 13188 21532 13198 21588
rect 34962 21532 34972 21588
rect 35028 21532 39340 21588
rect 39396 21532 42028 21588
rect 42084 21532 43484 21588
rect 43540 21532 43550 21588
rect 43652 21532 47628 21588
rect 47684 21532 47694 21588
rect 200 21504 800 21532
rect 43652 21476 43708 21532
rect 42914 21420 42924 21476
rect 42980 21420 43708 21476
rect 45042 21420 45052 21476
rect 45108 21420 45612 21476
rect 45668 21420 45678 21476
rect 51986 21196 51996 21252
rect 52052 21196 53676 21252
rect 53732 21196 53742 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 20850 20860 20860 20916
rect 20916 20860 24332 20916
rect 24388 20860 24398 20916
rect 24546 20860 24556 20916
rect 24612 20860 25340 20916
rect 25396 20860 25406 20916
rect 31154 20860 31164 20916
rect 31220 20860 32508 20916
rect 32564 20860 32574 20916
rect 45154 20748 45164 20804
rect 45220 20748 45948 20804
rect 46004 20748 46014 20804
rect 29810 20636 29820 20692
rect 29876 20636 30380 20692
rect 30436 20636 30446 20692
rect 2818 20524 2828 20580
rect 2884 20524 3836 20580
rect 3892 20524 3902 20580
rect 12338 20524 12348 20580
rect 12404 20524 13468 20580
rect 13524 20524 13534 20580
rect 35634 20524 35644 20580
rect 35700 20524 37548 20580
rect 37604 20524 37614 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 18722 20188 18732 20244
rect 18788 20188 19516 20244
rect 19572 20188 19582 20244
rect 26674 20188 26684 20244
rect 26740 20188 27468 20244
rect 27524 20188 27534 20244
rect 29698 20188 29708 20244
rect 29764 20188 32956 20244
rect 33012 20188 33022 20244
rect 33954 20188 33964 20244
rect 34020 20188 34860 20244
rect 34916 20188 37436 20244
rect 37492 20188 38108 20244
rect 38164 20188 38174 20244
rect 40002 20188 40012 20244
rect 40068 20188 40572 20244
rect 40628 20188 40638 20244
rect 49634 20188 49644 20244
rect 49700 20188 50540 20244
rect 50596 20188 50606 20244
rect 30604 20132 30660 20188
rect 30594 20076 30604 20132
rect 30660 20076 30670 20132
rect 36530 20076 36540 20132
rect 36596 20076 38444 20132
rect 38500 20076 38510 20132
rect 41458 20076 41468 20132
rect 41524 20076 42588 20132
rect 42644 20076 42654 20132
rect 43922 20076 43932 20132
rect 43988 20076 47180 20132
rect 47236 20076 47246 20132
rect 28802 19964 28812 20020
rect 28868 19964 30940 20020
rect 30996 19964 31006 20020
rect 36978 19964 36988 20020
rect 37044 19964 38332 20020
rect 38388 19964 38398 20020
rect 16818 19852 16828 19908
rect 16884 19852 18284 19908
rect 18340 19852 18350 19908
rect 22530 19852 22540 19908
rect 22596 19852 24556 19908
rect 24612 19852 25452 19908
rect 25508 19852 25518 19908
rect 37762 19852 37772 19908
rect 37828 19852 39340 19908
rect 39396 19852 39406 19908
rect 16930 19740 16940 19796
rect 16996 19740 17836 19796
rect 17892 19740 17902 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 5058 19404 5068 19460
rect 5124 19404 6300 19460
rect 6356 19404 6366 19460
rect 6738 19404 6748 19460
rect 6804 19404 8540 19460
rect 8596 19404 8606 19460
rect 4946 19292 4956 19348
rect 5012 19292 6076 19348
rect 6132 19292 6142 19348
rect 12562 19292 12572 19348
rect 12628 19292 13916 19348
rect 13972 19292 13982 19348
rect 15586 19292 15596 19348
rect 15652 19292 21532 19348
rect 21588 19292 21598 19348
rect 39890 19292 39900 19348
rect 39956 19292 40908 19348
rect 40964 19292 40974 19348
rect 38098 19180 38108 19236
rect 38164 19180 41356 19236
rect 41412 19180 41422 19236
rect 54898 19180 54908 19236
rect 54964 19180 56252 19236
rect 56308 19180 56812 19236
rect 56868 19180 56878 19236
rect 19170 19068 19180 19124
rect 19236 19068 19516 19124
rect 19572 19068 20076 19124
rect 20132 19068 22988 19124
rect 23044 19068 23054 19124
rect 52658 19068 52668 19124
rect 52724 19068 55580 19124
rect 55636 19068 55646 19124
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 19394 18508 19404 18564
rect 19460 18508 21196 18564
rect 21252 18508 22540 18564
rect 22596 18508 22764 18564
rect 22820 18508 22830 18564
rect 2146 18396 2156 18452
rect 2212 18396 7868 18452
rect 7924 18396 7934 18452
rect 14130 18396 14140 18452
rect 14196 18396 16436 18452
rect 16594 18396 16604 18452
rect 16660 18396 17948 18452
rect 18004 18396 19628 18452
rect 19684 18396 21308 18452
rect 21364 18396 21374 18452
rect 33394 18396 33404 18452
rect 33460 18396 40796 18452
rect 40852 18396 41916 18452
rect 41972 18396 41982 18452
rect 49634 18396 49644 18452
rect 49700 18396 51324 18452
rect 51380 18396 51390 18452
rect 16380 18340 16436 18396
rect 14802 18284 14812 18340
rect 14868 18284 15484 18340
rect 15540 18284 15550 18340
rect 16380 18284 17052 18340
rect 17108 18284 17276 18340
rect 17332 18284 17342 18340
rect 20738 18284 20748 18340
rect 20804 18284 21980 18340
rect 22036 18284 22046 18340
rect 33506 18284 33516 18340
rect 33572 18284 34636 18340
rect 34692 18284 34702 18340
rect 13122 18172 13132 18228
rect 13188 18172 17724 18228
rect 17780 18172 17790 18228
rect 22530 18172 22540 18228
rect 22596 18172 23324 18228
rect 23380 18172 23390 18228
rect 51762 18172 51772 18228
rect 51828 18172 53228 18228
rect 53284 18172 53294 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 13580 17836 19516 17892
rect 19572 17836 19582 17892
rect 13580 17780 13636 17836
rect 8372 17724 11788 17780
rect 11844 17724 13580 17780
rect 13636 17724 13646 17780
rect 46498 17724 46508 17780
rect 46564 17724 47628 17780
rect 47684 17724 47694 17780
rect 54786 17724 54796 17780
rect 54852 17724 55916 17780
rect 55972 17724 55982 17780
rect 8306 17612 8316 17668
rect 8372 17612 8428 17724
rect 41010 17500 41020 17556
rect 41076 17500 42364 17556
rect 42420 17500 42430 17556
rect 48290 17388 48300 17444
rect 48356 17388 48860 17444
rect 48916 17388 49644 17444
rect 49700 17388 49710 17444
rect 51986 17388 51996 17444
rect 52052 17388 52668 17444
rect 52724 17388 52734 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 25778 17052 25788 17108
rect 25844 17052 27580 17108
rect 27636 17052 28140 17108
rect 28196 17052 29036 17108
rect 29092 17052 29102 17108
rect 34738 17052 34748 17108
rect 34804 17052 37324 17108
rect 37380 17052 37390 17108
rect 47170 17052 47180 17108
rect 47236 17052 48748 17108
rect 48804 17052 49532 17108
rect 49588 17052 49598 17108
rect 32946 16940 32956 16996
rect 33012 16940 33740 16996
rect 33796 16940 33806 16996
rect 8978 16828 8988 16884
rect 9044 16828 9660 16884
rect 9716 16828 10780 16884
rect 10836 16828 11452 16884
rect 11508 16828 11518 16884
rect 19282 16828 19292 16884
rect 19348 16828 21756 16884
rect 21812 16828 21822 16884
rect 31042 16828 31052 16884
rect 31108 16828 33628 16884
rect 33684 16828 33694 16884
rect 36754 16828 36764 16884
rect 36820 16828 38556 16884
rect 38612 16828 38622 16884
rect 42802 16828 42812 16884
rect 42868 16828 45388 16884
rect 45444 16828 46060 16884
rect 46116 16828 46126 16884
rect 11452 16772 11508 16828
rect 5058 16716 5068 16772
rect 5124 16716 5740 16772
rect 5796 16716 8764 16772
rect 8820 16716 8830 16772
rect 11452 16716 12796 16772
rect 12852 16716 12862 16772
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 11554 16156 11564 16212
rect 11620 16156 13804 16212
rect 13860 16156 13870 16212
rect 37762 16156 37772 16212
rect 37828 16156 38780 16212
rect 38836 16156 38846 16212
rect 39778 16156 39788 16212
rect 39844 16156 40908 16212
rect 40964 16156 40974 16212
rect 44034 15932 44044 15988
rect 44100 15932 47628 15988
rect 47684 15932 47694 15988
rect 50530 15932 50540 15988
rect 50596 15932 53452 15988
rect 53508 15932 53518 15988
rect 22530 15820 22540 15876
rect 22596 15820 23772 15876
rect 23828 15820 23838 15876
rect 38882 15820 38892 15876
rect 38948 15820 41692 15876
rect 41748 15820 42140 15876
rect 42196 15820 44716 15876
rect 44772 15820 44782 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 49186 15372 49196 15428
rect 49252 15372 50316 15428
rect 50372 15372 50382 15428
rect 18834 15260 18844 15316
rect 18900 15260 19516 15316
rect 19572 15260 20412 15316
rect 20468 15260 20478 15316
rect 44482 15260 44492 15316
rect 44548 15260 45612 15316
rect 45668 15260 45678 15316
rect 13122 15148 13132 15204
rect 13188 15148 14364 15204
rect 14420 15148 14430 15204
rect 7970 15036 7980 15092
rect 8036 15036 8764 15092
rect 8820 15036 11340 15092
rect 11396 15036 11406 15092
rect 20178 15036 20188 15092
rect 20244 15036 20636 15092
rect 20692 15036 21420 15092
rect 21476 15036 21756 15092
rect 21812 15036 21822 15092
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 24658 14588 24668 14644
rect 24724 14588 27916 14644
rect 27972 14588 27982 14644
rect 39554 14588 39564 14644
rect 39620 14588 43820 14644
rect 43876 14588 46956 14644
rect 47012 14588 47022 14644
rect 50306 14588 50316 14644
rect 50372 14588 53116 14644
rect 53172 14588 53182 14644
rect 54114 14588 54124 14644
rect 54180 14588 55580 14644
rect 55636 14588 55646 14644
rect 16258 14252 16268 14308
rect 16324 14252 16828 14308
rect 16884 14252 17276 14308
rect 17332 14252 17342 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 21746 13916 21756 13972
rect 21812 13916 23884 13972
rect 23940 13916 23950 13972
rect 32050 13916 32060 13972
rect 32116 13916 33516 13972
rect 33572 13916 34076 13972
rect 34132 13916 35308 13972
rect 35364 13916 35374 13972
rect 8978 13804 8988 13860
rect 9044 13804 10500 13860
rect 10444 13748 10500 13804
rect 8642 13692 8652 13748
rect 8708 13692 9996 13748
rect 10052 13692 10062 13748
rect 10434 13692 10444 13748
rect 10500 13692 12572 13748
rect 12628 13692 12638 13748
rect 46946 13692 46956 13748
rect 47012 13692 47852 13748
rect 47908 13692 47918 13748
rect 52770 13692 52780 13748
rect 52836 13692 53564 13748
rect 53620 13692 53630 13748
rect 6290 13580 6300 13636
rect 6356 13580 6860 13636
rect 6916 13580 6926 13636
rect 25554 13468 25564 13524
rect 25620 13468 26236 13524
rect 26292 13468 29148 13524
rect 29204 13468 29214 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 16930 13132 16940 13188
rect 16996 13132 19292 13188
rect 19348 13132 19358 13188
rect 28466 13132 28476 13188
rect 28532 13132 29036 13188
rect 29092 13132 29102 13188
rect 4162 13020 4172 13076
rect 4228 13020 6972 13076
rect 7028 13020 7038 13076
rect 19954 13020 19964 13076
rect 20020 13020 23324 13076
rect 23380 13020 23390 13076
rect 41906 13020 41916 13076
rect 41972 13020 45836 13076
rect 45892 13020 45902 13076
rect 46274 13020 46284 13076
rect 46340 13020 47628 13076
rect 47684 13020 47694 13076
rect 6066 12908 6076 12964
rect 6132 12908 7308 12964
rect 7364 12908 7756 12964
rect 7812 12908 7822 12964
rect 8372 12908 8988 12964
rect 9044 12908 10668 12964
rect 10724 12908 10734 12964
rect 12562 12908 12572 12964
rect 12628 12908 13804 12964
rect 13860 12908 13870 12964
rect 35634 12908 35644 12964
rect 35700 12908 36316 12964
rect 36372 12908 36382 12964
rect 39106 12908 39116 12964
rect 39172 12908 41580 12964
rect 41636 12908 41646 12964
rect 8372 12852 8428 12908
rect 6850 12796 6860 12852
rect 6916 12796 8204 12852
rect 8260 12796 8428 12852
rect 9090 12796 9100 12852
rect 9156 12796 10332 12852
rect 10388 12796 10398 12852
rect 11330 12796 11340 12852
rect 11396 12796 11900 12852
rect 11956 12796 11966 12852
rect 14802 12796 14812 12852
rect 14868 12796 15596 12852
rect 15652 12796 15662 12852
rect 44034 12796 44044 12852
rect 44100 12796 46284 12852
rect 46340 12796 46350 12852
rect 4274 12684 4284 12740
rect 4340 12684 5740 12740
rect 5796 12684 6636 12740
rect 6692 12684 7756 12740
rect 7812 12684 7822 12740
rect 10994 12684 11004 12740
rect 11060 12684 11676 12740
rect 11732 12684 11742 12740
rect 13346 12684 13356 12740
rect 13412 12684 14028 12740
rect 14084 12684 14094 12740
rect 52210 12684 52220 12740
rect 52276 12684 53340 12740
rect 53396 12684 54460 12740
rect 54516 12684 54526 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 7186 12348 7196 12404
rect 7252 12348 9772 12404
rect 9828 12348 9838 12404
rect 33954 12348 33964 12404
rect 34020 12348 35532 12404
rect 35588 12348 35598 12404
rect 36978 12348 36988 12404
rect 37044 12348 38892 12404
rect 38948 12348 40236 12404
rect 40292 12348 40302 12404
rect 46386 12348 46396 12404
rect 46452 12348 48412 12404
rect 48468 12348 48478 12404
rect 53666 12348 53676 12404
rect 53732 12348 55020 12404
rect 55076 12348 56364 12404
rect 56420 12348 56430 12404
rect 8306 12124 8316 12180
rect 8372 12124 8988 12180
rect 9044 12124 9054 12180
rect 10994 12124 11004 12180
rect 11060 12124 13356 12180
rect 13412 12124 13422 12180
rect 13794 12124 13804 12180
rect 13860 12124 14476 12180
rect 14532 12124 14542 12180
rect 24098 12124 24108 12180
rect 24164 12124 28028 12180
rect 28084 12124 28094 12180
rect 41570 12124 41580 12180
rect 41636 12124 45276 12180
rect 45332 12124 45342 12180
rect 1922 12012 1932 12068
rect 1988 12012 3500 12068
rect 3556 12012 3948 12068
rect 4004 12012 5740 12068
rect 5796 12012 5806 12068
rect 9538 11900 9548 11956
rect 9604 11900 10108 11956
rect 10164 11900 11116 11956
rect 11172 11900 14252 11956
rect 14308 11900 14318 11956
rect 28354 11900 28364 11956
rect 28420 11900 32172 11956
rect 32228 11900 32238 11956
rect 12114 11788 12124 11844
rect 12180 11788 13020 11844
rect 13076 11788 15596 11844
rect 15652 11788 15662 11844
rect 29810 11788 29820 11844
rect 29876 11788 31948 11844
rect 32004 11788 32014 11844
rect 46050 11788 46060 11844
rect 46116 11788 46396 11844
rect 46452 11788 46462 11844
rect 54226 11788 54236 11844
rect 54292 11788 54302 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 54236 11732 54292 11788
rect 51986 11676 51996 11732
rect 52052 11676 54292 11732
rect 24994 11564 25004 11620
rect 25060 11564 25452 11620
rect 25508 11564 26124 11620
rect 26180 11564 26190 11620
rect 38322 11564 38332 11620
rect 38388 11564 38556 11620
rect 38612 11564 39116 11620
rect 39172 11564 40012 11620
rect 40068 11564 40078 11620
rect 44482 11564 44492 11620
rect 44548 11564 45724 11620
rect 45780 11564 45790 11620
rect 50754 11564 50764 11620
rect 50820 11564 53564 11620
rect 53620 11564 53630 11620
rect 16146 11452 16156 11508
rect 16212 11452 20412 11508
rect 20468 11452 26348 11508
rect 26404 11452 26414 11508
rect 35746 11452 35756 11508
rect 35812 11452 36204 11508
rect 36260 11452 39564 11508
rect 39620 11452 39630 11508
rect 50978 11452 50988 11508
rect 51044 11452 53676 11508
rect 53732 11452 53742 11508
rect 8194 11340 8204 11396
rect 8260 11340 10220 11396
rect 10276 11340 10286 11396
rect 47506 11340 47516 11396
rect 47572 11340 51996 11396
rect 52052 11340 52062 11396
rect 53442 11340 53452 11396
rect 53508 11340 54124 11396
rect 54180 11340 54190 11396
rect 6514 11228 6524 11284
rect 6580 11228 6748 11284
rect 6804 11228 6814 11284
rect 46386 11228 46396 11284
rect 46452 11228 47404 11284
rect 47460 11228 47470 11284
rect 10658 11116 10668 11172
rect 10724 11116 11004 11172
rect 11060 11116 11900 11172
rect 11956 11116 12236 11172
rect 12292 11116 12684 11172
rect 12740 11116 14028 11172
rect 14084 11116 14364 11172
rect 14420 11116 14430 11172
rect 38546 11116 38556 11172
rect 38612 11116 39228 11172
rect 39284 11116 39788 11172
rect 39844 11116 39854 11172
rect 45938 11116 45948 11172
rect 46004 11116 47180 11172
rect 47236 11116 47246 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 3154 10556 3164 10612
rect 3220 10556 4396 10612
rect 4452 10556 4462 10612
rect 7298 10556 7308 10612
rect 7364 10556 7374 10612
rect 8194 10556 8204 10612
rect 8260 10556 11004 10612
rect 11060 10556 11070 10612
rect 21970 10556 21980 10612
rect 22036 10556 22652 10612
rect 22708 10556 22718 10612
rect 50866 10556 50876 10612
rect 50932 10556 51436 10612
rect 51492 10556 51502 10612
rect 7308 10500 7364 10556
rect 2818 10444 2828 10500
rect 2884 10444 3948 10500
rect 4004 10444 4014 10500
rect 7308 10444 9772 10500
rect 9828 10444 9996 10500
rect 10052 10444 10062 10500
rect 22978 10444 22988 10500
rect 23044 10444 24668 10500
rect 24724 10444 24734 10500
rect 44706 10332 44716 10388
rect 44772 10332 45388 10388
rect 45444 10332 45454 10388
rect 19730 10220 19740 10276
rect 19796 10220 21868 10276
rect 21924 10220 21934 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 9874 10108 9884 10164
rect 9940 10108 11228 10164
rect 11284 10108 11294 10164
rect 38322 10108 38332 10164
rect 38388 10108 38780 10164
rect 38836 10108 38846 10164
rect 52434 10108 52444 10164
rect 52500 10108 53900 10164
rect 53956 10108 53966 10164
rect 45154 9996 45164 10052
rect 45220 9996 47852 10052
rect 47908 9996 48076 10052
rect 48132 9996 50876 10052
rect 50932 9996 50942 10052
rect 7186 9884 7196 9940
rect 7252 9884 8092 9940
rect 8148 9884 8158 9940
rect 16818 9884 16828 9940
rect 16884 9884 19068 9940
rect 19124 9884 19134 9940
rect 31938 9884 31948 9940
rect 32004 9884 33068 9940
rect 33124 9884 33134 9940
rect 39554 9884 39564 9940
rect 39620 9884 40460 9940
rect 40516 9884 40526 9940
rect 46610 9884 46620 9940
rect 46676 9884 47628 9940
rect 47684 9884 47694 9940
rect 54898 9884 54908 9940
rect 54964 9884 55580 9940
rect 55636 9884 55646 9940
rect 6962 9772 6972 9828
rect 7028 9772 8540 9828
rect 8596 9772 8606 9828
rect 12562 9772 12572 9828
rect 12628 9772 15596 9828
rect 15652 9772 15662 9828
rect 22194 9772 22204 9828
rect 22260 9772 22428 9828
rect 22484 9772 24668 9828
rect 24724 9772 24734 9828
rect 24882 9772 24892 9828
rect 24948 9772 27580 9828
rect 27636 9772 27646 9828
rect 4722 9660 4732 9716
rect 4788 9660 6748 9716
rect 6804 9660 7196 9716
rect 7252 9660 8316 9716
rect 8372 9660 8382 9716
rect 11330 9660 11340 9716
rect 11396 9660 11900 9716
rect 11956 9660 11966 9716
rect 7410 9548 7420 9604
rect 7476 9548 8652 9604
rect 8708 9548 8718 9604
rect 9314 9548 9324 9604
rect 9380 9548 10220 9604
rect 10276 9548 10780 9604
rect 10836 9548 10846 9604
rect 48626 9548 48636 9604
rect 48692 9548 50316 9604
rect 50372 9548 50382 9604
rect 6850 9436 6860 9492
rect 6916 9436 7868 9492
rect 7924 9436 7934 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 19058 9212 19068 9268
rect 19124 9212 20412 9268
rect 20468 9212 20478 9268
rect 24658 9212 24668 9268
rect 24724 9212 26908 9268
rect 26964 9212 26974 9268
rect 44594 9212 44604 9268
rect 44660 9212 45164 9268
rect 45220 9212 45230 9268
rect 3378 9100 3388 9156
rect 3444 9100 5964 9156
rect 6020 9100 6860 9156
rect 6916 9100 6926 9156
rect 7634 9100 7644 9156
rect 7700 9100 8876 9156
rect 8932 9100 8942 9156
rect 10994 9100 11004 9156
rect 11060 9100 13468 9156
rect 13524 9100 13534 9156
rect 4050 8988 4060 9044
rect 4116 8988 4732 9044
rect 4788 8988 4798 9044
rect 4946 8988 4956 9044
rect 5012 8988 6188 9044
rect 6244 8988 7420 9044
rect 7476 8988 7486 9044
rect 7970 8988 7980 9044
rect 8036 8988 8540 9044
rect 8596 8988 8606 9044
rect 12786 8988 12796 9044
rect 12852 8988 13356 9044
rect 13412 8988 15484 9044
rect 15540 8988 15708 9044
rect 15764 8988 16044 9044
rect 16100 8988 16828 9044
rect 16884 8988 16894 9044
rect 37650 8988 37660 9044
rect 37716 8988 40236 9044
rect 40292 8988 40684 9044
rect 40740 8988 41020 9044
rect 41076 8988 41804 9044
rect 41860 8988 41870 9044
rect 41804 8932 41860 8988
rect 41804 8876 44380 8932
rect 44436 8876 44446 8932
rect 8978 8764 8988 8820
rect 9044 8764 10220 8820
rect 10276 8764 10286 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 22082 8428 22092 8484
rect 22148 8428 22876 8484
rect 22932 8428 22942 8484
rect 6514 8316 6524 8372
rect 6580 8316 10108 8372
rect 10164 8316 10174 8372
rect 49074 8316 49084 8372
rect 49140 8316 51324 8372
rect 51380 8316 51772 8372
rect 51828 8316 52668 8372
rect 52724 8316 52734 8372
rect 20850 8204 20860 8260
rect 20916 8204 21868 8260
rect 21924 8204 24444 8260
rect 24500 8204 24510 8260
rect 48738 8204 48748 8260
rect 48804 8204 49756 8260
rect 49812 8204 49822 8260
rect 51874 8204 51884 8260
rect 51940 8204 54124 8260
rect 54180 8204 54190 8260
rect 10098 8092 10108 8148
rect 10164 8092 11004 8148
rect 11060 8092 11070 8148
rect 19618 7980 19628 8036
rect 19684 7980 20748 8036
rect 20804 7980 20814 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 29922 7644 29932 7700
rect 29988 7644 30492 7700
rect 30548 7644 30558 7700
rect 55234 7644 55244 7700
rect 55300 7644 55692 7700
rect 55748 7644 56252 7700
rect 56308 7644 56318 7700
rect 2146 7532 2156 7588
rect 2212 7532 3948 7588
rect 4004 7532 4844 7588
rect 4900 7532 5740 7588
rect 5796 7532 8540 7588
rect 8596 7532 8606 7588
rect 12114 7532 12124 7588
rect 12180 7532 14700 7588
rect 14756 7532 14766 7588
rect 24658 7532 24668 7588
rect 24724 7532 26236 7588
rect 26292 7532 27804 7588
rect 27860 7532 27870 7588
rect 43250 7532 43260 7588
rect 43316 7532 45500 7588
rect 45556 7532 45566 7588
rect 54450 7532 54460 7588
rect 54516 7532 55356 7588
rect 55412 7532 55422 7588
rect 2594 7420 2604 7476
rect 2660 7420 3724 7476
rect 3780 7420 3790 7476
rect 20626 7420 20636 7476
rect 20692 7420 22092 7476
rect 22148 7420 23100 7476
rect 23156 7420 23166 7476
rect 26562 7420 26572 7476
rect 26628 7420 27132 7476
rect 27188 7420 27916 7476
rect 27972 7420 27982 7476
rect 38210 7420 38220 7476
rect 38276 7420 38780 7476
rect 38836 7420 39228 7476
rect 39284 7420 39294 7476
rect 10770 7308 10780 7364
rect 10836 7308 11452 7364
rect 11508 7308 12012 7364
rect 12068 7308 12078 7364
rect 19954 7308 19964 7364
rect 20020 7308 22652 7364
rect 22708 7308 22718 7364
rect 27794 7308 27804 7364
rect 27860 7308 29260 7364
rect 29316 7308 29326 7364
rect 38546 7308 38556 7364
rect 38612 7308 39116 7364
rect 39172 7308 39182 7364
rect 52322 7308 52332 7364
rect 52388 7308 53564 7364
rect 53620 7308 53630 7364
rect 22754 7196 22764 7252
rect 22820 7196 24444 7252
rect 24500 7196 25564 7252
rect 25620 7196 26796 7252
rect 26852 7196 27356 7252
rect 27412 7196 27422 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 52546 6860 52556 6916
rect 52612 6860 53788 6916
rect 53844 6860 53854 6916
rect 11330 6748 11340 6804
rect 11396 6748 12236 6804
rect 12292 6748 12302 6804
rect 46274 6748 46284 6804
rect 46340 6748 48972 6804
rect 49028 6748 49420 6804
rect 49476 6748 49644 6804
rect 49700 6748 49710 6804
rect 52658 6748 52668 6804
rect 52724 6748 53340 6804
rect 53396 6748 53406 6804
rect 11900 6692 11956 6748
rect 2258 6636 2268 6692
rect 2324 6636 2716 6692
rect 2772 6636 4172 6692
rect 4228 6636 4238 6692
rect 11890 6636 11900 6692
rect 11956 6636 11966 6692
rect 15810 6636 15820 6692
rect 15876 6636 19180 6692
rect 19236 6636 22092 6692
rect 22148 6636 22158 6692
rect 26562 6636 26572 6692
rect 26628 6636 27244 6692
rect 27300 6636 27310 6692
rect 39778 6636 39788 6692
rect 39844 6636 40012 6692
rect 40068 6636 40460 6692
rect 40516 6636 40526 6692
rect 49074 6636 49084 6692
rect 49140 6636 54012 6692
rect 54068 6636 54078 6692
rect 3714 6524 3724 6580
rect 3780 6524 9100 6580
rect 9156 6524 9166 6580
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 22082 6076 22092 6132
rect 22148 6076 22428 6132
rect 22484 6076 23212 6132
rect 23268 6076 23660 6132
rect 23716 6076 26236 6132
rect 26292 6076 26302 6132
rect 2818 5964 2828 6020
rect 2884 5964 3948 6020
rect 4004 5964 4014 6020
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 59200 5460 59800 5488
rect 55346 5404 55356 5460
rect 55412 5404 59800 5460
rect 59200 5376 59800 5404
rect 40114 5180 40124 5236
rect 40180 5180 41244 5236
rect 41300 5180 41310 5236
rect 40562 5068 40572 5124
rect 40628 5068 40908 5124
rect 40964 5068 41916 5124
rect 41972 5068 43932 5124
rect 43988 5068 43998 5124
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 18 3612 28 3668
rect 84 3612 2492 3668
rect 2548 3612 2558 3668
rect 21522 3612 21532 3668
rect 21588 3612 22428 3668
rect 22484 3612 22494 3668
rect 43698 3612 43708 3668
rect 43764 3612 45612 3668
rect 45668 3612 45678 3668
rect 43362 3500 43372 3556
rect 43428 3500 44940 3556
rect 44996 3500 45006 3556
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0493__A2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 49616 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0503__A4
timestamp 1669390400
transform 1 0 36736 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0504__A2
timestamp 1669390400
transform 1 0 39200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0513__I
timestamp 1669390400
transform 1 0 8960 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0543__A2
timestamp 1669390400
transform 1 0 9072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0561__A3
timestamp 1669390400
transform 1 0 50400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0572__I
timestamp 1669390400
transform -1 0 2352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0586__A1
timestamp 1669390400
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0589__A1
timestamp 1669390400
transform 1 0 9632 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0595__A2
timestamp 1669390400
transform 1 0 25536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0598__A2
timestamp 1669390400
transform -1 0 26880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0600__A1
timestamp 1669390400
transform 1 0 26096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0607__A1
timestamp 1669390400
transform -1 0 22736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0630__A1
timestamp 1669390400
transform 1 0 9408 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0631__A2
timestamp 1669390400
transform 1 0 39088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0633__A1
timestamp 1669390400
transform 1 0 39984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0636__A1
timestamp 1669390400
transform 1 0 38752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0644__A3
timestamp 1669390400
transform 1 0 14000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0648__A1
timestamp 1669390400
transform -1 0 4256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0648__A2
timestamp 1669390400
transform -1 0 3808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0650__A1
timestamp 1669390400
transform 1 0 4368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0650__A2
timestamp 1669390400
transform 1 0 3920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0656__I
timestamp 1669390400
transform 1 0 10640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0660__A2
timestamp 1669390400
transform 1 0 10976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0663__A1
timestamp 1669390400
transform 1 0 12768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0665__A2
timestamp 1669390400
transform 1 0 9296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0666__A2
timestamp 1669390400
transform 1 0 11872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0671__B2
timestamp 1669390400
transform 1 0 7728 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0676__B
timestamp 1669390400
transform 1 0 47488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0697__A2
timestamp 1669390400
transform -1 0 48944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0705__I
timestamp 1669390400
transform 1 0 26880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0706__A2
timestamp 1669390400
transform 1 0 29456 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0708__A1
timestamp 1669390400
transform 1 0 27776 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0711__A2
timestamp 1669390400
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0714__A2
timestamp 1669390400
transform -1 0 29008 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0716__A1
timestamp 1669390400
transform -1 0 26656 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0719__A2
timestamp 1669390400
transform 1 0 26656 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0723__B
timestamp 1669390400
transform -1 0 27216 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0725__CLK
timestamp 1669390400
transform 1 0 17024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0726__CLK
timestamp 1669390400
transform 1 0 16352 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0727__CLK
timestamp 1669390400
transform 1 0 12880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0728__CLK
timestamp 1669390400
transform 1 0 8064 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0731__CLK
timestamp 1669390400
transform 1 0 5600 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0732__CLK
timestamp 1669390400
transform 1 0 4368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0733__CLK
timestamp 1669390400
transform -1 0 18928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0734__CLK
timestamp 1669390400
transform -1 0 17248 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0735__CLK
timestamp 1669390400
transform 1 0 13552 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0736__CLK
timestamp 1669390400
transform 1 0 11648 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0737__CLK
timestamp 1669390400
transform 1 0 17584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0738__CLK
timestamp 1669390400
transform 1 0 16576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0739__CLK
timestamp 1669390400
transform 1 0 12432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0740__CLK
timestamp 1669390400
transform 1 0 11200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0741__CLK
timestamp 1669390400
transform 1 0 7728 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0742__CLK
timestamp 1669390400
transform 1 0 8736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__CLK
timestamp 1669390400
transform 1 0 12432 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0744__CLK
timestamp 1669390400
transform -1 0 9856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0745__CLK
timestamp 1669390400
transform 1 0 12320 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0746__CLK
timestamp 1669390400
transform 1 0 10864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0747__CLK
timestamp 1669390400
transform -1 0 8176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0748__CLK
timestamp 1669390400
transform 1 0 9296 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0749__CLK
timestamp 1669390400
transform 1 0 5824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0750__CLK
timestamp 1669390400
transform 1 0 4928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0751__CLK
timestamp 1669390400
transform -1 0 5824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0752__CLK
timestamp 1669390400
transform 1 0 53312 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0752__D
timestamp 1669390400
transform 1 0 56896 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0753__CLK
timestamp 1669390400
transform 1 0 26208 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0754__CLK
timestamp 1669390400
transform 1 0 30464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0756__CLK
timestamp 1669390400
transform 1 0 23632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0757__CLK
timestamp 1669390400
transform 1 0 23296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0758__CLK
timestamp 1669390400
transform 1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0759__CLK
timestamp 1669390400
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0760__CLK
timestamp 1669390400
transform 1 0 21280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0761__CLK
timestamp 1669390400
transform 1 0 20608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0762__CLK
timestamp 1669390400
transform 1 0 25536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0763__CLK
timestamp 1669390400
transform -1 0 21392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0764__CLK
timestamp 1669390400
transform 1 0 19824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0765__CLK
timestamp 1669390400
transform 1 0 22624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0766__CLK
timestamp 1669390400
transform 1 0 25760 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0768__CLK
timestamp 1669390400
transform 1 0 20160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0769__CLK
timestamp 1669390400
transform 1 0 29008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0772__CLK
timestamp 1669390400
transform 1 0 33040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0773__CLK
timestamp 1669390400
transform 1 0 33488 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__CLK
timestamp 1669390400
transform 1 0 36736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0775__CLK
timestamp 1669390400
transform 1 0 16240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0776__CLK
timestamp 1669390400
transform 1 0 17248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__CLK
timestamp 1669390400
transform 1 0 19040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0778__CLK
timestamp 1669390400
transform 1 0 19152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__CLK
timestamp 1669390400
transform -1 0 23520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0780__CLK
timestamp 1669390400
transform 1 0 23856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0781__CLK
timestamp 1669390400
transform 1 0 4928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0782__CLK
timestamp 1669390400
transform 1 0 54096 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__CLK
timestamp 1669390400
transform 1 0 52304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0785__CLK
timestamp 1669390400
transform 1 0 45472 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0787__CLK
timestamp 1669390400
transform -1 0 37632 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__CLK
timestamp 1669390400
transform 1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0789__CLK
timestamp 1669390400
transform 1 0 36064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0790__CLK
timestamp 1669390400
transform 1 0 35168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0791__CLK
timestamp 1669390400
transform 1 0 33264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0792__CLK
timestamp 1669390400
transform 1 0 39424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0794__CLK
timestamp 1669390400
transform 1 0 34720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0795__CLK
timestamp 1669390400
transform 1 0 38080 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0796__CLK
timestamp 1669390400
transform 1 0 36960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0797__CLK
timestamp 1669390400
transform 1 0 31584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0798__CLK
timestamp 1669390400
transform 1 0 32928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0799__CLK
timestamp 1669390400
transform 1 0 31920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0800__CLK
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0801__CLK
timestamp 1669390400
transform 1 0 41440 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0803__CLK
timestamp 1669390400
transform 1 0 46144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0805__CLK
timestamp 1669390400
transform -1 0 42448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0806__CLK
timestamp 1669390400
transform 1 0 41440 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0807__CLK
timestamp 1669390400
transform 1 0 43792 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0808__CLK
timestamp 1669390400
transform 1 0 45360 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0809__CLK
timestamp 1669390400
transform -1 0 35392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0810__CLK
timestamp 1669390400
transform -1 0 44016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0811__CLK
timestamp 1669390400
transform 1 0 9632 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0812__CLK
timestamp 1669390400
transform 1 0 6384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0813__CLK
timestamp 1669390400
transform -1 0 6944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0814__CLK
timestamp 1669390400
transform 1 0 11200 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0815__CLK
timestamp 1669390400
transform 1 0 21616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0816__CLK
timestamp 1669390400
transform -1 0 27888 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0817__CLK
timestamp 1669390400
transform 1 0 27328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0818__CLK
timestamp 1669390400
transform 1 0 29568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0819__CLK
timestamp 1669390400
transform 1 0 25536 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0820__CLK
timestamp 1669390400
transform -1 0 21840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0821__CLK
timestamp 1669390400
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0822__CLK
timestamp 1669390400
transform 1 0 28112 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0823__CLK
timestamp 1669390400
transform 1 0 19376 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0824__CLK
timestamp 1669390400
transform 1 0 20832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0825__CLK
timestamp 1669390400
transform 1 0 21616 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0826__CLK
timestamp 1669390400
transform -1 0 20160 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__CLK
timestamp 1669390400
transform 1 0 20832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0828__CLK
timestamp 1669390400
transform 1 0 18256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__CLK
timestamp 1669390400
transform 1 0 22176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0830__CLK
timestamp 1669390400
transform -1 0 21056 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0831__CLK
timestamp 1669390400
transform 1 0 13104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0832__CLK
timestamp 1669390400
transform 1 0 13552 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__CLK
timestamp 1669390400
transform 1 0 16576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0834__CLK
timestamp 1669390400
transform -1 0 16464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0835__CLK
timestamp 1669390400
transform -1 0 17248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__CLK
timestamp 1669390400
transform 1 0 12208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0837__CLK
timestamp 1669390400
transform 1 0 16128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0838__CLK
timestamp 1669390400
transform 1 0 18256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0839__CLK
timestamp 1669390400
transform 1 0 48944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0840__CLK
timestamp 1669390400
transform 1 0 40208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0841__CLK
timestamp 1669390400
transform 1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__CLK
timestamp 1669390400
transform 1 0 40880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0843__CLK
timestamp 1669390400
transform 1 0 38864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0844__CLK
timestamp 1669390400
transform 1 0 42112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0845__CLK
timestamp 1669390400
transform 1 0 38080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0846__CLK
timestamp 1669390400
transform 1 0 37408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0847__CLK
timestamp 1669390400
transform 1 0 41328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__CLK
timestamp 1669390400
transform 1 0 38528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0849__CLK
timestamp 1669390400
transform 1 0 34048 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__CLK
timestamp 1669390400
transform 1 0 27552 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__CLK
timestamp 1669390400
transform 1 0 33936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0852__CLK
timestamp 1669390400
transform 1 0 35280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0853__CLK
timestamp 1669390400
transform 1 0 35056 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0855__CLK
timestamp 1669390400
transform 1 0 34720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0857__CLK
timestamp 1669390400
transform 1 0 30464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__CLK
timestamp 1669390400
transform 1 0 32704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__CLK
timestamp 1669390400
transform 1 0 31808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__CLK
timestamp 1669390400
transform 1 0 32256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__CLK
timestamp 1669390400
transform -1 0 28112 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0865__CLK
timestamp 1669390400
transform 1 0 32928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__CLK
timestamp 1669390400
transform 1 0 38752 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0868__CLK
timestamp 1669390400
transform 1 0 52752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__CLK
timestamp 1669390400
transform 1 0 46368 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__CLK
timestamp 1669390400
transform 1 0 47152 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__CLK
timestamp 1669390400
transform 1 0 50512 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__CLK
timestamp 1669390400
transform 1 0 52640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__CLK
timestamp 1669390400
transform -1 0 53088 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__CLK
timestamp 1669390400
transform 1 0 54208 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__CLK
timestamp 1669390400
transform 1 0 53312 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0876__CLK
timestamp 1669390400
transform 1 0 52640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__CLK
timestamp 1669390400
transform 1 0 54544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0878__CLK
timestamp 1669390400
transform 1 0 56336 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__CLK
timestamp 1669390400
transform 1 0 47040 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__CLK
timestamp 1669390400
transform 1 0 44688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__CLK
timestamp 1669390400
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0882__CLK
timestamp 1669390400
transform -1 0 49056 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0886__CLK
timestamp 1669390400
transform 1 0 44912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0887__CLK
timestamp 1669390400
transform -1 0 40880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0888__CLK
timestamp 1669390400
transform 1 0 38528 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__CLK
timestamp 1669390400
transform 1 0 44352 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__CLK
timestamp 1669390400
transform 1 0 36736 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0891__CLK
timestamp 1669390400
transform -1 0 37520 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__CLK
timestamp 1669390400
transform 1 0 36960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__CLK
timestamp 1669390400
transform -1 0 37184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__CLK
timestamp 1669390400
transform 1 0 36288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0895__CLK
timestamp 1669390400
transform 1 0 41440 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__CLK
timestamp 1669390400
transform 1 0 39424 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0898__CLK
timestamp 1669390400
transform 1 0 54992 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__CLK
timestamp 1669390400
transform 1 0 51408 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0902__CLK
timestamp 1669390400
transform 1 0 48832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__CLK
timestamp 1669390400
transform 1 0 44352 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__CLK
timestamp 1669390400
transform 1 0 40208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__CLK
timestamp 1669390400
transform 1 0 41888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__CLK
timestamp 1669390400
transform 1 0 48832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__CLK
timestamp 1669390400
transform 1 0 48272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__CLK
timestamp 1669390400
transform 1 0 44688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__CLK
timestamp 1669390400
transform 1 0 46032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__CLK
timestamp 1669390400
transform 1 0 48832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0911__CLK
timestamp 1669390400
transform 1 0 53312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__CLK
timestamp 1669390400
transform 1 0 50736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0913__CLK
timestamp 1669390400
transform 1 0 52864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0914__CLK
timestamp 1669390400
transform 1 0 56784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__CLK
timestamp 1669390400
transform 1 0 51968 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0916__CLK
timestamp 1669390400
transform 1 0 52640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0917__CLK
timestamp 1669390400
transform 1 0 56784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0918__CLK
timestamp 1669390400
transform 1 0 57120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__CLK
timestamp 1669390400
transform 1 0 51744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0920__CLK
timestamp 1669390400
transform 1 0 49392 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__CLK
timestamp 1669390400
transform 1 0 53312 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0922__CLK
timestamp 1669390400
transform 1 0 55664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__CLK
timestamp 1669390400
transform 1 0 52640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__CLK
timestamp 1669390400
transform 1 0 56784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0926__CLK
timestamp 1669390400
transform -1 0 53312 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__CLK
timestamp 1669390400
transform 1 0 15904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0933__CLK
timestamp 1669390400
transform 1 0 16016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__CLK
timestamp 1669390400
transform 1 0 14000 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0935__CLK
timestamp 1669390400
transform -1 0 11424 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0937__CLK
timestamp 1669390400
transform 1 0 12768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0938__CLK
timestamp 1669390400
transform 1 0 13552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__CLK
timestamp 1669390400
transform 1 0 10752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__CLK
timestamp 1669390400
transform -1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__CLK
timestamp 1669390400
transform 1 0 9632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0942__CLK
timestamp 1669390400
transform 1 0 13104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__CLK
timestamp 1669390400
transform 1 0 12320 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0944__CLK
timestamp 1669390400
transform 1 0 11984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0945__CLK
timestamp 1669390400
transform 1 0 13552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0946__CLK
timestamp 1669390400
transform 1 0 17024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0947__CLK
timestamp 1669390400
transform 1 0 14112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0948__CLK
timestamp 1669390400
transform -1 0 17360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0949__CLK
timestamp 1669390400
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__CLK
timestamp 1669390400
transform 1 0 5712 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0951__CLK
timestamp 1669390400
transform 1 0 5600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0952__CLK
timestamp 1669390400
transform -1 0 5376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__CLK
timestamp 1669390400
transform 1 0 5600 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0954__CLK
timestamp 1669390400
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__CLK
timestamp 1669390400
transform 1 0 27664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0956__CLK
timestamp 1669390400
transform 1 0 44912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0957__CLK
timestamp 1669390400
transform 1 0 46816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0958__CLK
timestamp 1669390400
transform 1 0 45360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0959__CLK
timestamp 1669390400
transform 1 0 48496 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0960__CLK
timestamp 1669390400
transform 1 0 51296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__CLK
timestamp 1669390400
transform 1 0 54880 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0962__CLK
timestamp 1669390400
transform -1 0 56000 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0963__CLK
timestamp 1669390400
transform 1 0 53312 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0964__CLK
timestamp 1669390400
transform 1 0 48048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0965__CLK
timestamp 1669390400
transform 1 0 42336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0966__CLK
timestamp 1669390400
transform 1 0 42560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__CLK
timestamp 1669390400
transform 1 0 36960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0969__CLK
timestamp 1669390400
transform 1 0 40432 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0970__CLK
timestamp 1669390400
transform 1 0 40880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__CLK
timestamp 1669390400
transform 1 0 43344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0975__CLK
timestamp 1669390400
transform 1 0 44912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__CLK
timestamp 1669390400
transform 1 0 40768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0977__CLK
timestamp 1669390400
transform 1 0 46144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0978__CLK
timestamp 1669390400
transform 1 0 46704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0979__CLK
timestamp 1669390400
transform 1 0 45696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__CLK
timestamp 1669390400
transform 1 0 41440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__CLK
timestamp 1669390400
transform 1 0 31696 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__CLK
timestamp 1669390400
transform 1 0 30912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__CLK
timestamp 1669390400
transform 1 0 34160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__CLK
timestamp 1669390400
transform 1 0 31136 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0990__CLK
timestamp 1669390400
transform 1 0 20832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0991__CLK
timestamp 1669390400
transform 1 0 28112 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0992__CLK
timestamp 1669390400
transform -1 0 26320 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0993__CLK
timestamp 1669390400
transform 1 0 21504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0994__CLK
timestamp 1669390400
transform 1 0 20832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__CLK
timestamp 1669390400
transform 1 0 23520 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0996__CLK
timestamp 1669390400
transform 1 0 22736 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0997__CLK
timestamp 1669390400
transform 1 0 27888 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__CLK
timestamp 1669390400
transform 1 0 27888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1000__CLK
timestamp 1669390400
transform -1 0 25760 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__CLK
timestamp 1669390400
transform -1 0 17808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1002__CLK
timestamp 1669390400
transform 1 0 21056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__CLK
timestamp 1669390400
transform 1 0 24416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1004__CLK
timestamp 1669390400
transform 1 0 22960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1005__CLK
timestamp 1669390400
transform 1 0 23296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1006__CLK
timestamp 1669390400
transform -1 0 22064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__CLK
timestamp 1669390400
transform 1 0 17584 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1008__CLK
timestamp 1669390400
transform 1 0 20944 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__CLK
timestamp 1669390400
transform 1 0 22848 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__CLK
timestamp 1669390400
transform 1 0 17584 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1011__CLK
timestamp 1669390400
transform 1 0 21616 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__CLK
timestamp 1669390400
transform 1 0 23184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1013__CLK
timestamp 1669390400
transform 1 0 22400 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1014__CLK
timestamp 1669390400
transform -1 0 13328 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1669390400
transform -1 0 28336 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clk_I
timestamp 1669390400
transform 1 0 21504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clk_I
timestamp 1669390400
transform 1 0 18704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clk_I
timestamp 1669390400
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clk_I
timestamp 1669390400
transform -1 0 41440 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_0_clk_I
timestamp 1669390400
transform 1 0 9184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_1_clk_I
timestamp 1669390400
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_2_clk_I
timestamp 1669390400
transform 1 0 11200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_3_clk_I
timestamp 1669390400
transform 1 0 17024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_4_clk_I
timestamp 1669390400
transform 1 0 23408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_5_clk_I
timestamp 1669390400
transform -1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_6_clk_I
timestamp 1669390400
transform 1 0 18480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_7_clk_I
timestamp 1669390400
transform 1 0 13664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_8_clk_I
timestamp 1669390400
transform -1 0 15456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_9_clk_I
timestamp 1669390400
transform 1 0 12656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_10_clk_I
timestamp 1669390400
transform 1 0 15792 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_11_clk_I
timestamp 1669390400
transform 1 0 10752 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_12_clk_I
timestamp 1669390400
transform -1 0 9856 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_13_clk_I
timestamp 1669390400
transform 1 0 13552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_14_clk_I
timestamp 1669390400
transform 1 0 16912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_15_clk_I
timestamp 1669390400
transform 1 0 26432 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_16_clk_I
timestamp 1669390400
transform 1 0 26656 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_17_clk_I
timestamp 1669390400
transform 1 0 19040 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_18_clk_I
timestamp 1669390400
transform 1 0 24192 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_19_clk_I
timestamp 1669390400
transform 1 0 36736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_20_clk_I
timestamp 1669390400
transform 1 0 39984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_21_clk_I
timestamp 1669390400
transform 1 0 44352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_22_clk_I
timestamp 1669390400
transform 1 0 40208 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_23_clk_I
timestamp 1669390400
transform -1 0 42336 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_24_clk_I
timestamp 1669390400
transform 1 0 49392 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_25_clk_I
timestamp 1669390400
transform 1 0 48720 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_26_clk_I
timestamp 1669390400
transform 1 0 50848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_27_clk_I
timestamp 1669390400
transform 1 0 46816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_29_clk_I
timestamp 1669390400
transform 1 0 46816 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_30_clk_I
timestamp 1669390400
transform 1 0 48048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_31_clk_I
timestamp 1669390400
transform -1 0 44240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_32_clk_I
timestamp 1669390400
transform 1 0 42784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_33_clk_I
timestamp 1669390400
transform 1 0 47264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_34_clk_I
timestamp 1669390400
transform -1 0 49392 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_35_clk_I
timestamp 1669390400
transform 1 0 50848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_36_clk_I
timestamp 1669390400
transform 1 0 48720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_37_clk_I
timestamp 1669390400
transform 1 0 50848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_38_clk_I
timestamp 1669390400
transform 1 0 48048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_39_clk_I
timestamp 1669390400
transform 1 0 47824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_40_clk_I
timestamp 1669390400
transform 1 0 45136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_41_clk_I
timestamp 1669390400
transform 1 0 36176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_42_clk_I
timestamp 1669390400
transform 1 0 43792 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_43_clk_I
timestamp 1669390400
transform 1 0 39312 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_44_clk_I
timestamp 1669390400
transform 1 0 26320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_45_clk_I
timestamp 1669390400
transform 1 0 22960 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_46_clk_I
timestamp 1669390400
transform 1 0 18816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_47_clk_I
timestamp 1669390400
transform 1 0 26320 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_48_clk_I
timestamp 1669390400
transform 1 0 19040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_49_clk_I
timestamp 1669390400
transform 1 0 20384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_50_clk_I
timestamp 1669390400
transform 1 0 9184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output8_I
timestamp 1669390400
transform -1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5040 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5488 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1669390400
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_177 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_195 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23184 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_203
timestamp 1669390400
transform 1 0 24080 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_207
timestamp 1669390400
transform 1 0 24528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1669390400
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_402
timestamp 1669390400
transform 1 0 46368 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_418
timestamp 1669390400
transform 1 0 48160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1669390400
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1669390400
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_508
timestamp 1669390400
transform 1 0 58240 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1669390400
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1669390400
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1669390400
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1669390400
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1669390400
transform 1 0 40544 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_421
timestamp 1669390400
transform 1 0 48496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1669390400
transform 1 0 56448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1669390400
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_507
timestamp 1669390400
transform 1 0 58128 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1669390400
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1669390400
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1669390400
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1669390400
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_337
timestamp 1669390400
transform 1 0 39088 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_345
timestamp 1669390400
transform 1 0 39984 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_347
timestamp 1669390400
transform 1 0 40208 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_377
timestamp 1669390400
transform 1 0 43568 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_381
timestamp 1669390400
transform 1 0 44016 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_456
timestamp 1669390400
transform 1 0 52416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1669390400
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_471
timestamp 1669390400
transform 1 0 54096 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_475
timestamp 1669390400
transform 1 0 54544 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_491
timestamp 1669390400
transform 1 0 56336 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_507
timestamp 1669390400
transform 1 0 58128 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_32
timestamp 1669390400
transform 1 0 4928 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_64
timestamp 1669390400
transform 1 0 8512 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_68
timestamp 1669390400
transform 1 0 8960 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_89
timestamp 1669390400
transform 1 0 11312 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_98
timestamp 1669390400
transform 1 0 12320 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_130
timestamp 1669390400
transform 1 0 15904 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_138
timestamp 1669390400
transform 1 0 16800 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_152
timestamp 1669390400
transform 1 0 18368 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_156
timestamp 1669390400
transform 1 0 18816 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_186
timestamp 1669390400
transform 1 0 22176 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_190
timestamp 1669390400
transform 1 0 22624 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_206
timestamp 1669390400
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_210
timestamp 1669390400
transform 1 0 24864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_219
timestamp 1669390400
transform 1 0 25872 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_221
timestamp 1669390400
transform 1 0 26096 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_224
timestamp 1669390400
transform 1 0 26432 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_256
timestamp 1669390400
transform 1 0 30016 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_272
timestamp 1669390400
transform 1 0 31808 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_280
timestamp 1669390400
transform 1 0 32704 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_318
timestamp 1669390400
transform 1 0 36960 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_334
timestamp 1669390400
transform 1 0 38752 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_340
timestamp 1669390400
transform 1 0 39424 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_348
timestamp 1669390400
transform 1 0 40320 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_352
timestamp 1669390400
transform 1 0 40768 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1669390400
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_431
timestamp 1669390400
transform 1 0 49616 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_447
timestamp 1669390400
transform 1 0 51408 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_455
timestamp 1669390400
transform 1 0 52304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_461
timestamp 1669390400
transform 1 0 52976 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1669390400
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1669390400
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_507
timestamp 1669390400
transform 1 0 58128 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_6
timestamp 1669390400
transform 1 0 2016 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_9
timestamp 1669390400
transform 1 0 2352 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_15
timestamp 1669390400
transform 1 0 3024 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_19
timestamp 1669390400
transform 1 0 3472 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_22
timestamp 1669390400
transform 1 0 3808 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_26
timestamp 1669390400
transform 1 0 4256 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_53
timestamp 1669390400
transform 1 0 7280 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_61
timestamp 1669390400
transform 1 0 8176 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_91
timestamp 1669390400
transform 1 0 11536 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1669390400
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1669390400
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_183
timestamp 1669390400
transform 1 0 21840 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_187
timestamp 1669390400
transform 1 0 22288 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_191
timestamp 1669390400
transform 1 0 22736 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_222
timestamp 1669390400
transform 1 0 26208 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_228
timestamp 1669390400
transform 1 0 26880 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_238
timestamp 1669390400
transform 1 0 28000 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_246
timestamp 1669390400
transform 1 0 28896 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_351
timestamp 1669390400
transform 1 0 40656 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_355
timestamp 1669390400
transform 1 0 41104 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_387
timestamp 1669390400
transform 1 0 44688 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_396
timestamp 1669390400
transform 1 0 45696 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_398
timestamp 1669390400
transform 1 0 45920 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_428
timestamp 1669390400
transform 1 0 49280 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_459
timestamp 1669390400
transform 1 0 52752 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_466
timestamp 1669390400
transform 1 0 53536 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_498
timestamp 1669390400
transform 1 0 57120 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_506
timestamp 1669390400
transform 1 0 58016 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_508
timestamp 1669390400
transform 1 0 58240 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_18
timestamp 1669390400
transform 1 0 3360 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_75
timestamp 1669390400
transform 1 0 9744 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_89
timestamp 1669390400
transform 1 0 11312 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_97
timestamp 1669390400
transform 1 0 12208 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_128
timestamp 1669390400
transform 1 0 15680 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_132
timestamp 1669390400
transform 1 0 16128 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_140
timestamp 1669390400
transform 1 0 17024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_152
timestamp 1669390400
transform 1 0 18368 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_156
timestamp 1669390400
transform 1 0 18816 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_187
timestamp 1669390400
transform 1 0 22288 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_195
timestamp 1669390400
transform 1 0 23184 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_201
timestamp 1669390400
transform 1 0 23856 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_211
timestamp 1669390400
transform 1 0 24976 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_218
timestamp 1669390400
transform 1 0 25760 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_220
timestamp 1669390400
transform 1 0 25984 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_227
timestamp 1669390400
transform 1 0 26768 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_258
timestamp 1669390400
transform 1 0 30240 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_262
timestamp 1669390400
transform 1 0 30688 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_278
timestamp 1669390400
transform 1 0 32480 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_282
timestamp 1669390400
transform 1 0 32928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_318
timestamp 1669390400
transform 1 0 36960 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_326
timestamp 1669390400
transform 1 0 37856 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_334
timestamp 1669390400
transform 1 0 38752 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_348
timestamp 1669390400
transform 1 0 40320 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_352
timestamp 1669390400
transform 1 0 40768 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_361
timestamp 1669390400
transform 1 0 41776 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_364
timestamp 1669390400
transform 1 0 42112 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_395
timestamp 1669390400
transform 1 0 45584 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_411
timestamp 1669390400
transform 1 0 47376 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_419
timestamp 1669390400
transform 1 0 48272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_423
timestamp 1669390400
transform 1 0 48720 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_440
timestamp 1669390400
transform 1 0 50624 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_448
timestamp 1669390400
transform 1 0 51520 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_452
timestamp 1669390400
transform 1 0 51968 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_483
timestamp 1669390400
transform 1 0 55440 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_487
timestamp 1669390400
transform 1 0 55888 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_495
timestamp 1669390400
transform 1 0 56784 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_507
timestamp 1669390400
transform 1 0 58128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_4
timestamp 1669390400
transform 1 0 1792 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_67
timestamp 1669390400
transform 1 0 8848 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_69
timestamp 1669390400
transform 1 0 9072 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_72
timestamp 1669390400
transform 1 0 9408 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_82
timestamp 1669390400
transform 1 0 10528 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_97
timestamp 1669390400
transform 1 0 12208 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_124
timestamp 1669390400
transform 1 0 15232 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_157
timestamp 1669390400
transform 1 0 18928 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_161
timestamp 1669390400
transform 1 0 19376 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_169
timestamp 1669390400
transform 1 0 20272 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_189
timestamp 1669390400
transform 1 0 22512 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_197
timestamp 1669390400
transform 1 0 23408 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_230
timestamp 1669390400
transform 1 0 27104 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_240
timestamp 1669390400
transform 1 0 28224 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_329
timestamp 1669390400
transform 1 0 38192 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_333
timestamp 1669390400
transform 1 0 38640 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_336
timestamp 1669390400
transform 1 0 38976 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_338
timestamp 1669390400
transform 1 0 39200 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_397
timestamp 1669390400
transform 1 0 45808 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_405
timestamp 1669390400
transform 1 0 46704 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_407
timestamp 1669390400
transform 1 0 46928 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_412
timestamp 1669390400
transform 1 0 47488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_420
timestamp 1669390400
transform 1 0 48384 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_453
timestamp 1669390400
transform 1 0 52080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_457
timestamp 1669390400
transform 1 0 52528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_474
timestamp 1669390400
transform 1 0 54432 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_506
timestamp 1669390400
transform 1 0 58016 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_508
timestamp 1669390400
transform 1 0 58240 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_10
timestamp 1669390400
transform 1 0 2464 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_14
timestamp 1669390400
transform 1 0 2912 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_28
timestamp 1669390400
transform 1 0 4480 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_36
timestamp 1669390400
transform 1 0 5376 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_46
timestamp 1669390400
transform 1 0 6496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_50
timestamp 1669390400
transform 1 0 6944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_62
timestamp 1669390400
transform 1 0 8288 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_84
timestamp 1669390400
transform 1 0 10752 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_88
timestamp 1669390400
transform 1 0 11200 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_96
timestamp 1669390400
transform 1 0 12096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_129
timestamp 1669390400
transform 1 0 15792 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_133
timestamp 1669390400
transform 1 0 16240 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_152
timestamp 1669390400
transform 1 0 18368 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_156
timestamp 1669390400
transform 1 0 18816 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_160
timestamp 1669390400
transform 1 0 19264 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_223
timestamp 1669390400
transform 1 0 26320 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_227
timestamp 1669390400
transform 1 0 26768 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_239
timestamp 1669390400
transform 1 0 28112 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_255
timestamp 1669390400
transform 1 0 29904 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_259
timestamp 1669390400
transform 1 0 30352 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_265
timestamp 1669390400
transform 1 0 31024 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_281
timestamp 1669390400
transform 1 0 32816 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_318
timestamp 1669390400
transform 1 0 36960 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_326
timestamp 1669390400
transform 1 0 37856 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_330
timestamp 1669390400
transform 1 0 38304 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_344
timestamp 1669390400
transform 1 0 39872 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_346
timestamp 1669390400
transform 1 0 40096 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_349
timestamp 1669390400
transform 1 0 40432 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_353
timestamp 1669390400
transform 1 0 40880 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_359
timestamp 1669390400
transform 1 0 41552 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_389
timestamp 1669390400
transform 1 0 44912 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_393
timestamp 1669390400
transform 1 0 45360 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_409
timestamp 1669390400
transform 1 0 47152 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_419
timestamp 1669390400
transform 1 0 48272 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_479
timestamp 1669390400
transform 1 0 54992 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_485
timestamp 1669390400
transform 1 0 55664 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_493
timestamp 1669390400
transform 1 0 56560 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_507
timestamp 1669390400
transform 1 0 58128 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_32
timestamp 1669390400
transform 1 0 4928 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_45
timestamp 1669390400
transform 1 0 6384 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_56
timestamp 1669390400
transform 1 0 7616 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_66
timestamp 1669390400
transform 1 0 8736 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_70
timestamp 1669390400
transform 1 0 9184 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_73
timestamp 1669390400
transform 1 0 9520 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_81
timestamp 1669390400
transform 1 0 10416 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_91
timestamp 1669390400
transform 1 0 11536 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_124
timestamp 1669390400
transform 1 0 15232 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_126
timestamp 1669390400
transform 1 0 15456 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_156
timestamp 1669390400
transform 1 0 18816 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_160
timestamp 1669390400
transform 1 0 19264 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_191
timestamp 1669390400
transform 1 0 22736 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_199
timestamp 1669390400
transform 1 0 23632 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_203
timestamp 1669390400
transform 1 0 24080 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_212
timestamp 1669390400
transform 1 0 25088 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_228
timestamp 1669390400
transform 1 0 26880 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_237
timestamp 1669390400
transform 1 0 27888 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_245
timestamp 1669390400
transform 1 0 28784 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_281
timestamp 1669390400
transform 1 0 32816 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_285
timestamp 1669390400
transform 1 0 33264 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_317
timestamp 1669390400
transform 1 0 36848 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_351
timestamp 1669390400
transform 1 0 40656 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_382
timestamp 1669390400
transform 1 0 44128 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_386
timestamp 1669390400
transform 1 0 44576 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_422
timestamp 1669390400
transform 1 0 48608 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_426
timestamp 1669390400
transform 1 0 49056 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_428
timestamp 1669390400
transform 1 0 49280 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_458
timestamp 1669390400
transform 1 0 52640 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_493
timestamp 1669390400
transform 1 0 56560 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_497
timestamp 1669390400
transform 1 0 57008 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_505
timestamp 1669390400
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_10
timestamp 1669390400
transform 1 0 2464 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_12
timestamp 1669390400
transform 1 0 2688 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_21
timestamp 1669390400
transform 1 0 3696 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_25
timestamp 1669390400
transform 1 0 4144 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_29
timestamp 1669390400
transform 1 0 4592 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_45
timestamp 1669390400
transform 1 0 6384 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_56
timestamp 1669390400
transform 1 0 7616 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_64
timestamp 1669390400
transform 1 0 8512 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_68
timestamp 1669390400
transform 1 0 8960 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_80
timestamp 1669390400
transform 1 0 10304 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_88
timestamp 1669390400
transform 1 0 11200 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_92
timestamp 1669390400
transform 1 0 11648 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_94
timestamp 1669390400
transform 1 0 11872 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_100
timestamp 1669390400
transform 1 0 12544 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_104
timestamp 1669390400
transform 1 0 12992 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_140
timestamp 1669390400
transform 1 0 17024 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_152
timestamp 1669390400
transform 1 0 18368 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_185
timestamp 1669390400
transform 1 0 22064 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_194
timestamp 1669390400
transform 1 0 23072 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_198
timestamp 1669390400
transform 1 0 23520 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_206
timestamp 1669390400
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_210
timestamp 1669390400
transform 1 0 24864 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_223
timestamp 1669390400
transform 1 0 26320 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_227
timestamp 1669390400
transform 1 0 26768 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_241
timestamp 1669390400
transform 1 0 28336 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_318
timestamp 1669390400
transform 1 0 36960 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_326
timestamp 1669390400
transform 1 0 37856 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_336
timestamp 1669390400
transform 1 0 38976 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_343
timestamp 1669390400
transform 1 0 39760 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_347
timestamp 1669390400
transform 1 0 40208 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_363
timestamp 1669390400
transform 1 0 42000 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_367
timestamp 1669390400
transform 1 0 42448 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_373
timestamp 1669390400
transform 1 0 43120 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_389
timestamp 1669390400
transform 1 0 44912 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_400
timestamp 1669390400
transform 1 0 46144 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_406
timestamp 1669390400
transform 1 0 46816 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_414
timestamp 1669390400
transform 1 0 47712 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_418
timestamp 1669390400
transform 1 0 48160 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_424
timestamp 1669390400
transform 1 0 48832 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_436
timestamp 1669390400
transform 1 0 50176 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_440
timestamp 1669390400
transform 1 0 50624 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_444
timestamp 1669390400
transform 1 0 51072 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_507
timestamp 1669390400
transform 1 0 58128 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_67
timestamp 1669390400
transform 1 0 8848 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_69
timestamp 1669390400
transform 1 0 9072 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_72
timestamp 1669390400
transform 1 0 9408 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_74
timestamp 1669390400
transform 1 0 9632 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_81
timestamp 1669390400
transform 1 0 10416 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_85
timestamp 1669390400
transform 1 0 10864 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_93
timestamp 1669390400
transform 1 0 11760 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_96
timestamp 1669390400
transform 1 0 12096 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_112
timestamp 1669390400
transform 1 0 13888 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_115
timestamp 1669390400
transform 1 0 14224 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_117
timestamp 1669390400
transform 1 0 14448 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_168
timestamp 1669390400
transform 1 0 20160 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_189
timestamp 1669390400
transform 1 0 22512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_193
timestamp 1669390400
transform 1 0 22960 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_195
timestamp 1669390400
transform 1 0 23184 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_212
timestamp 1669390400
transform 1 0 25088 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_258
timestamp 1669390400
transform 1 0 30240 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_309
timestamp 1669390400
transform 1 0 35952 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_313
timestamp 1669390400
transform 1 0 36400 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_317
timestamp 1669390400
transform 1 0 36848 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_335
timestamp 1669390400
transform 1 0 38864 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_339
timestamp 1669390400
transform 1 0 39312 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_371
timestamp 1669390400
transform 1 0 42896 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_387
timestamp 1669390400
transform 1 0 44688 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_404
timestamp 1669390400
transform 1 0 46592 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_413
timestamp 1669390400
transform 1 0 47600 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_415
timestamp 1669390400
transform 1 0 47824 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_445
timestamp 1669390400
transform 1 0 51184 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_449
timestamp 1669390400
transform 1 0 51632 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_457
timestamp 1669390400
transform 1 0 52528 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_474
timestamp 1669390400
transform 1 0 54432 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_480
timestamp 1669390400
transform 1 0 55104 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_496
timestamp 1669390400
transform 1 0 56896 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_504
timestamp 1669390400
transform 1 0 57792 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_508
timestamp 1669390400
transform 1 0 58240 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_18
timestamp 1669390400
transform 1 0 3360 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_82
timestamp 1669390400
transform 1 0 10528 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_113
timestamp 1669390400
transform 1 0 14000 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_131
timestamp 1669390400
transform 1 0 16016 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_139
timestamp 1669390400
transform 1 0 16912 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_160
timestamp 1669390400
transform 1 0 19264 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_164
timestamp 1669390400
transform 1 0 19712 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_194
timestamp 1669390400
transform 1 0 23072 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_198
timestamp 1669390400
transform 1 0 23520 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_207
timestamp 1669390400
transform 1 0 24528 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_211
timestamp 1669390400
transform 1 0 24976 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_219
timestamp 1669390400
transform 1 0 25872 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_223
timestamp 1669390400
transform 1 0 26320 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_231
timestamp 1669390400
transform 1 0 27216 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_235
timestamp 1669390400
transform 1 0 27664 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_245
timestamp 1669390400
transform 1 0 28784 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_276
timestamp 1669390400
transform 1 0 32256 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_288
timestamp 1669390400
transform 1 0 33600 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_293
timestamp 1669390400
transform 1 0 34160 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_309
timestamp 1669390400
transform 1 0 35952 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_313
timestamp 1669390400
transform 1 0 36400 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_315
timestamp 1669390400
transform 1 0 36624 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_345
timestamp 1669390400
transform 1 0 39984 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_349
timestamp 1669390400
transform 1 0 40432 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_353
timestamp 1669390400
transform 1 0 40880 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_387
timestamp 1669390400
transform 1 0 44688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_391
timestamp 1669390400
transform 1 0 45136 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_422
timestamp 1669390400
transform 1 0 48608 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_433
timestamp 1669390400
transform 1 0 49840 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_437
timestamp 1669390400
transform 1 0 50288 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_439
timestamp 1669390400
transform 1 0 50512 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_469
timestamp 1669390400
transform 1 0 53872 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_477
timestamp 1669390400
transform 1 0 54768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_481
timestamp 1669390400
transform 1 0 55216 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_507
timestamp 1669390400
transform 1 0 58128 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_44
timestamp 1669390400
transform 1 0 6272 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_55
timestamp 1669390400
transform 1 0 7504 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_59
timestamp 1669390400
transform 1 0 7952 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_63
timestamp 1669390400
transform 1 0 8400 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_65
timestamp 1669390400
transform 1 0 8624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_74
timestamp 1669390400
transform 1 0 9632 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_82
timestamp 1669390400
transform 1 0 10528 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_91
timestamp 1669390400
transform 1 0 11536 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_112
timestamp 1669390400
transform 1 0 13888 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_115
timestamp 1669390400
transform 1 0 14224 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_123
timestamp 1669390400
transform 1 0 15120 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_125
timestamp 1669390400
transform 1 0 15344 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_130
timestamp 1669390400
transform 1 0 15904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_134
timestamp 1669390400
transform 1 0 16352 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_140
timestamp 1669390400
transform 1 0 17024 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_144
timestamp 1669390400
transform 1 0 17472 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_152
timestamp 1669390400
transform 1 0 18368 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_154
timestamp 1669390400
transform 1 0 18592 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_167
timestamp 1669390400
transform 1 0 20048 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_175
timestamp 1669390400
transform 1 0 20944 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_184
timestamp 1669390400
transform 1 0 21952 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_206
timestamp 1669390400
transform 1 0 24416 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_222
timestamp 1669390400
transform 1 0 26208 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_225
timestamp 1669390400
transform 1 0 26544 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_233
timestamp 1669390400
transform 1 0 27440 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_245
timestamp 1669390400
transform 1 0 28784 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_283
timestamp 1669390400
transform 1 0 33040 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_329
timestamp 1669390400
transform 1 0 38192 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_333
timestamp 1669390400
transform 1 0 38640 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_364
timestamp 1669390400
transform 1 0 42112 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_372
timestamp 1669390400
transform 1 0 43008 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_376
timestamp 1669390400
transform 1 0 43456 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_378
timestamp 1669390400
transform 1 0 43680 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_383
timestamp 1669390400
transform 1 0 44240 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_387
timestamp 1669390400
transform 1 0 44688 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_422
timestamp 1669390400
transform 1 0 48608 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_426
timestamp 1669390400
transform 1 0 49056 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_458
timestamp 1669390400
transform 1 0 52640 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_473
timestamp 1669390400
transform 1 0 54320 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_505
timestamp 1669390400
transform 1 0 57904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_10
timestamp 1669390400
transform 1 0 2464 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_14
timestamp 1669390400
transform 1 0 2912 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_16
timestamp 1669390400
transform 1 0 3136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_46
timestamp 1669390400
transform 1 0 6496 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_52
timestamp 1669390400
transform 1 0 7168 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_56
timestamp 1669390400
transform 1 0 7616 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_92
timestamp 1669390400
transform 1 0 11648 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_108
timestamp 1669390400
transform 1 0 13440 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_150
timestamp 1669390400
transform 1 0 18144 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_166
timestamp 1669390400
transform 1 0 19936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_199
timestamp 1669390400
transform 1 0 23632 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_203
timestamp 1669390400
transform 1 0 24080 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_211
timestamp 1669390400
transform 1 0 24976 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_223
timestamp 1669390400
transform 1 0 26320 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_275
timestamp 1669390400
transform 1 0 32144 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_289
timestamp 1669390400
transform 1 0 33712 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_297
timestamp 1669390400
transform 1 0 34608 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_301
timestamp 1669390400
transform 1 0 35056 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_332
timestamp 1669390400
transform 1 0 38528 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_336
timestamp 1669390400
transform 1 0 38976 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_348
timestamp 1669390400
transform 1 0 40320 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_352
timestamp 1669390400
transform 1 0 40768 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_361
timestamp 1669390400
transform 1 0 41776 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_413
timestamp 1669390400
transform 1 0 47600 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_417
timestamp 1669390400
transform 1 0 48048 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_460
timestamp 1669390400
transform 1 0 52864 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_471
timestamp 1669390400
transform 1 0 54096 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_487
timestamp 1669390400
transform 1 0 55888 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_495
timestamp 1669390400
transform 1 0 56784 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_507
timestamp 1669390400
transform 1 0 58128 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_53
timestamp 1669390400
transform 1 0 7280 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_86
timestamp 1669390400
transform 1 0 10976 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_90
timestamp 1669390400
transform 1 0 11424 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_124
timestamp 1669390400
transform 1 0 15232 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_132
timestamp 1669390400
transform 1 0 16128 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_135
timestamp 1669390400
transform 1 0 16464 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_166
timestamp 1669390400
transform 1 0 19936 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_170
timestamp 1669390400
transform 1 0 20384 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_210
timestamp 1669390400
transform 1 0 24864 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_241
timestamp 1669390400
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_245
timestamp 1669390400
transform 1 0 28784 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_254
timestamp 1669390400
transform 1 0 29792 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_259
timestamp 1669390400
transform 1 0 30352 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_267
timestamp 1669390400
transform 1 0 31248 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_271
timestamp 1669390400
transform 1 0 31696 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_301
timestamp 1669390400
transform 1 0 35056 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_305
timestamp 1669390400
transform 1 0 35504 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_309
timestamp 1669390400
transform 1 0 35952 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_315
timestamp 1669390400
transform 1 0 36624 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_325
timestamp 1669390400
transform 1 0 37744 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_377
timestamp 1669390400
transform 1 0 43568 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_381
timestamp 1669390400
transform 1 0 44016 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_396
timestamp 1669390400
transform 1 0 45696 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_398
timestamp 1669390400
transform 1 0 45920 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_403
timestamp 1669390400
transform 1 0 46480 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_407
timestamp 1669390400
transform 1 0 46928 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_409
timestamp 1669390400
transform 1 0 47152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_439
timestamp 1669390400
transform 1 0 50512 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_443
timestamp 1669390400
transform 1 0 50960 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_459
timestamp 1669390400
transform 1 0 52752 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_493
timestamp 1669390400
transform 1 0 56560 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_497
timestamp 1669390400
transform 1 0 57008 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_505
timestamp 1669390400
transform 1 0 57904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_75
timestamp 1669390400
transform 1 0 9744 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_80
timestamp 1669390400
transform 1 0 10304 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_96
timestamp 1669390400
transform 1 0 12096 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_133
timestamp 1669390400
transform 1 0 16240 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_152
timestamp 1669390400
transform 1 0 18368 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_158
timestamp 1669390400
transform 1 0 19040 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_210
timestamp 1669390400
transform 1 0 24864 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_219
timestamp 1669390400
transform 1 0 25872 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_249
timestamp 1669390400
transform 1 0 29232 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_281
timestamp 1669390400
transform 1 0 32816 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_302
timestamp 1669390400
transform 1 0 35168 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_333
timestamp 1669390400
transform 1 0 38640 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_337
timestamp 1669390400
transform 1 0 39088 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_353
timestamp 1669390400
transform 1 0 40880 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_361
timestamp 1669390400
transform 1 0 41776 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_367
timestamp 1669390400
transform 1 0 42448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_383
timestamp 1669390400
transform 1 0 44240 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_391
timestamp 1669390400
transform 1 0 45136 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_393
timestamp 1669390400
transform 1 0 45360 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_404
timestamp 1669390400
transform 1 0 46592 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_412
timestamp 1669390400
transform 1 0 47488 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_416
timestamp 1669390400
transform 1 0 47936 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_418
timestamp 1669390400
transform 1 0 48160 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_423
timestamp 1669390400
transform 1 0 48720 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_458
timestamp 1669390400
transform 1 0 52640 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_462
timestamp 1669390400
transform 1 0 53088 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_466
timestamp 1669390400
transform 1 0 53536 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_468
timestamp 1669390400
transform 1 0 53760 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_473
timestamp 1669390400
transform 1 0 54320 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_489
timestamp 1669390400
transform 1 0 56112 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_507
timestamp 1669390400
transform 1 0 58128 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_18
timestamp 1669390400
transform 1 0 3360 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_26
timestamp 1669390400
transform 1 0 4256 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_31
timestamp 1669390400
transform 1 0 4816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_40
timestamp 1669390400
transform 1 0 5824 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_56
timestamp 1669390400
transform 1 0 7616 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_93
timestamp 1669390400
transform 1 0 11760 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_95
timestamp 1669390400
transform 1 0 11984 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_100
timestamp 1669390400
transform 1 0 12544 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_104
timestamp 1669390400
transform 1 0 12992 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_119
timestamp 1669390400
transform 1 0 14672 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_127
timestamp 1669390400
transform 1 0 15568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_131
timestamp 1669390400
transform 1 0 16016 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_133
timestamp 1669390400
transform 1 0 16240 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_163
timestamp 1669390400
transform 1 0 19600 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_167
timestamp 1669390400
transform 1 0 20048 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_175
timestamp 1669390400
transform 1 0 20944 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_195
timestamp 1669390400
transform 1 0 23184 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_203
timestamp 1669390400
transform 1 0 24080 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_219
timestamp 1669390400
transform 1 0 25872 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_227
timestamp 1669390400
transform 1 0 26768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_233
timestamp 1669390400
transform 1 0 27440 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_241
timestamp 1669390400
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_245
timestamp 1669390400
transform 1 0 28784 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_254
timestamp 1669390400
transform 1 0 29792 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_284
timestamp 1669390400
transform 1 0 33152 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_290
timestamp 1669390400
transform 1 0 33824 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_294
timestamp 1669390400
transform 1 0 34272 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_310
timestamp 1669390400
transform 1 0 36064 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_316
timestamp 1669390400
transform 1 0 36736 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_331
timestamp 1669390400
transform 1 0 38416 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_362
timestamp 1669390400
transform 1 0 41888 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_366
timestamp 1669390400
transform 1 0 42336 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_374
timestamp 1669390400
transform 1 0 43232 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_378
timestamp 1669390400
transform 1 0 43680 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_383
timestamp 1669390400
transform 1 0 44240 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_422
timestamp 1669390400
transform 1 0 48608 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_424
timestamp 1669390400
transform 1 0 48832 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_429
timestamp 1669390400
transform 1 0 49392 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_468
timestamp 1669390400
transform 1 0 53760 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_500
timestamp 1669390400
transform 1 0 57344 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_508
timestamp 1669390400
transform 1 0 58240 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_35
timestamp 1669390400
transform 1 0 5264 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_78
timestamp 1669390400
transform 1 0 10080 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_82
timestamp 1669390400
transform 1 0 10528 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_86
timestamp 1669390400
transform 1 0 10976 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_117
timestamp 1669390400
transform 1 0 14448 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_123
timestamp 1669390400
transform 1 0 15120 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_139
timestamp 1669390400
transform 1 0 16912 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_149
timestamp 1669390400
transform 1 0 18032 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_157
timestamp 1669390400
transform 1 0 18928 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_188
timestamp 1669390400
transform 1 0 22400 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_192
timestamp 1669390400
transform 1 0 22848 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_194
timestamp 1669390400
transform 1 0 23072 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_203
timestamp 1669390400
transform 1 0 24080 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_211
timestamp 1669390400
transform 1 0 24976 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_217
timestamp 1669390400
transform 1 0 25648 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_220
timestamp 1669390400
transform 1 0 25984 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_228
timestamp 1669390400
transform 1 0 26880 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_232
timestamp 1669390400
transform 1 0 27328 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_236
timestamp 1669390400
transform 1 0 27776 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_267
timestamp 1669390400
transform 1 0 31248 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_273
timestamp 1669390400
transform 1 0 31920 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_281
timestamp 1669390400
transform 1 0 32816 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_305
timestamp 1669390400
transform 1 0 35504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_313
timestamp 1669390400
transform 1 0 36400 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_315
timestamp 1669390400
transform 1 0 36624 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_318
timestamp 1669390400
transform 1 0 36960 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_336
timestamp 1669390400
transform 1 0 38976 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_340
timestamp 1669390400
transform 1 0 39424 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_345
timestamp 1669390400
transform 1 0 39984 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_353
timestamp 1669390400
transform 1 0 40880 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_365
timestamp 1669390400
transform 1 0 42224 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_367
timestamp 1669390400
transform 1 0 42448 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_397
timestamp 1669390400
transform 1 0 45808 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_401
timestamp 1669390400
transform 1 0 46256 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_417
timestamp 1669390400
transform 1 0 48048 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_479
timestamp 1669390400
transform 1 0 54992 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_495
timestamp 1669390400
transform 1 0 56784 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_507
timestamp 1669390400
transform 1 0 58128 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_49
timestamp 1669390400
transform 1 0 6832 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_53
timestamp 1669390400
transform 1 0 7280 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_111
timestamp 1669390400
transform 1 0 13776 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_127
timestamp 1669390400
transform 1 0 15568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_135
timestamp 1669390400
transform 1 0 16464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_139
timestamp 1669390400
transform 1 0 16912 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_143
timestamp 1669390400
transform 1 0 17360 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_151
timestamp 1669390400
transform 1 0 18256 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_159
timestamp 1669390400
transform 1 0 19152 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_171
timestamp 1669390400
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_175
timestamp 1669390400
transform 1 0 20944 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_187
timestamp 1669390400
transform 1 0 22288 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_218
timestamp 1669390400
transform 1 0 25760 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_222
timestamp 1669390400
transform 1 0 26208 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_227
timestamp 1669390400
transform 1 0 26768 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1669390400
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_255
timestamp 1669390400
transform 1 0 29904 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_287
timestamp 1669390400
transform 1 0 33488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_295
timestamp 1669390400
transform 1 0 34384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_299
timestamp 1669390400
transform 1 0 34832 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_304
timestamp 1669390400
transform 1 0 35392 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_312
timestamp 1669390400
transform 1 0 36288 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_316
timestamp 1669390400
transform 1 0 36736 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_337
timestamp 1669390400
transform 1 0 39088 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_345
timestamp 1669390400
transform 1 0 39984 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_349
timestamp 1669390400
transform 1 0 40432 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_351
timestamp 1669390400
transform 1 0 40656 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_356
timestamp 1669390400
transform 1 0 41216 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_387
timestamp 1669390400
transform 1 0 44688 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_422
timestamp 1669390400
transform 1 0 48608 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_426
timestamp 1669390400
transform 1 0 49056 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_442
timestamp 1669390400
transform 1 0 50848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_450
timestamp 1669390400
transform 1 0 51744 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_454
timestamp 1669390400
transform 1 0 52192 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_496
timestamp 1669390400
transform 1 0 56896 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_500
timestamp 1669390400
transform 1 0 57344 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_508
timestamp 1669390400
transform 1 0 58240 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_36
timestamp 1669390400
transform 1 0 5376 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_52
timestamp 1669390400
transform 1 0 7168 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_68
timestamp 1669390400
transform 1 0 8960 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_81
timestamp 1669390400
transform 1 0 10416 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_86
timestamp 1669390400
transform 1 0 10976 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_94
timestamp 1669390400
transform 1 0 11872 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_98
timestamp 1669390400
transform 1 0 12320 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_110
timestamp 1669390400
transform 1 0 13664 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_175
timestamp 1669390400
transform 1 0 20944 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_179
timestamp 1669390400
transform 1 0 21392 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_191
timestamp 1669390400
transform 1 0 22736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_195
timestamp 1669390400
transform 1 0 23184 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_201
timestamp 1669390400
transform 1 0 23856 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_209
timestamp 1669390400
transform 1 0 24752 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_245
timestamp 1669390400
transform 1 0 28784 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_249
timestamp 1669390400
transform 1 0 29232 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_265
timestamp 1669390400
transform 1 0 31024 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_273
timestamp 1669390400
transform 1 0 31920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_281
timestamp 1669390400
transform 1 0 32816 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_290
timestamp 1669390400
transform 1 0 33824 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_320
timestamp 1669390400
transform 1 0 37184 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_324
timestamp 1669390400
transform 1 0 37632 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_332
timestamp 1669390400
transform 1 0 38528 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_338
timestamp 1669390400
transform 1 0 39200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_346
timestamp 1669390400
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_411
timestamp 1669390400
transform 1 0 47376 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_419
timestamp 1669390400
transform 1 0 48272 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_423
timestamp 1669390400
transform 1 0 48720 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_458
timestamp 1669390400
transform 1 0 52640 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_460
timestamp 1669390400
transform 1 0 52864 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_471
timestamp 1669390400
transform 1 0 54096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_479
timestamp 1669390400
transform 1 0 54992 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_495
timestamp 1669390400
transform 1 0 56784 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_507
timestamp 1669390400
transform 1 0 58128 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_4
timestamp 1669390400
transform 1 0 1792 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_53
timestamp 1669390400
transform 1 0 7280 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_69
timestamp 1669390400
transform 1 0 9072 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_102
timestamp 1669390400
transform 1 0 12768 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_111
timestamp 1669390400
transform 1 0 13776 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_119
timestamp 1669390400
transform 1 0 14672 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_123
timestamp 1669390400
transform 1 0 15120 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_174
timestamp 1669390400
transform 1 0 20832 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_182
timestamp 1669390400
transform 1 0 21728 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_190
timestamp 1669390400
transform 1 0 22624 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_192
timestamp 1669390400
transform 1 0 22848 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_195
timestamp 1669390400
transform 1 0 23184 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_258
timestamp 1669390400
transform 1 0 30240 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_289
timestamp 1669390400
transform 1 0 33712 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_293
timestamp 1669390400
transform 1 0 34160 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_309
timestamp 1669390400
transform 1 0 35952 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_317
timestamp 1669390400
transform 1 0 36848 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_325
timestamp 1669390400
transform 1 0 37744 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_355
timestamp 1669390400
transform 1 0 41104 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_359
timestamp 1669390400
transform 1 0 41552 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_375
timestamp 1669390400
transform 1 0 43344 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_383
timestamp 1669390400
transform 1 0 44240 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_387
timestamp 1669390400
transform 1 0 44688 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_400
timestamp 1669390400
transform 1 0 46144 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_405
timestamp 1669390400
transform 1 0 46704 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_421
timestamp 1669390400
transform 1 0 48496 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_452
timestamp 1669390400
transform 1 0 51968 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_493
timestamp 1669390400
transform 1 0 56560 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_497
timestamp 1669390400
transform 1 0 57008 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_505
timestamp 1669390400
transform 1 0 57904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_35
timestamp 1669390400
transform 1 0 5264 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_79
timestamp 1669390400
transform 1 0 10192 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_81
timestamp 1669390400
transform 1 0 10416 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_86
timestamp 1669390400
transform 1 0 10976 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_102
timestamp 1669390400
transform 1 0 12768 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_110
timestamp 1669390400
transform 1 0 13664 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_140
timestamp 1669390400
transform 1 0 17024 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_155
timestamp 1669390400
transform 1 0 18704 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_159
timestamp 1669390400
transform 1 0 19152 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_165
timestamp 1669390400
transform 1 0 19824 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_169
timestamp 1669390400
transform 1 0 20272 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_171
timestamp 1669390400
transform 1 0 20496 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_174
timestamp 1669390400
transform 1 0 20832 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_205
timestamp 1669390400
transform 1 0 24304 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_209
timestamp 1669390400
transform 1 0 24752 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_218
timestamp 1669390400
transform 1 0 25760 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_226
timestamp 1669390400
transform 1 0 26656 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_230
timestamp 1669390400
transform 1 0 27104 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_236
timestamp 1669390400
transform 1 0 27776 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_256
timestamp 1669390400
transform 1 0 30016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_260
timestamp 1669390400
transform 1 0 30464 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_262
timestamp 1669390400
transform 1 0 30688 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_269
timestamp 1669390400
transform 1 0 31472 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_277
timestamp 1669390400
transform 1 0 32368 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_281
timestamp 1669390400
transform 1 0 32816 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_290
timestamp 1669390400
transform 1 0 33824 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_296
timestamp 1669390400
transform 1 0 34496 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_327
timestamp 1669390400
transform 1 0 37968 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_347
timestamp 1669390400
transform 1 0 40208 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_353
timestamp 1669390400
transform 1 0 40880 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_373
timestamp 1669390400
transform 1 0 43120 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_381
timestamp 1669390400
transform 1 0 44016 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_389
timestamp 1669390400
transform 1 0 44912 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_419
timestamp 1669390400
transform 1 0 48272 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_423
timestamp 1669390400
transform 1 0 48720 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_436
timestamp 1669390400
transform 1 0 50176 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_442
timestamp 1669390400
transform 1 0 50848 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_446
timestamp 1669390400
transform 1 0 51296 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_476
timestamp 1669390400
transform 1 0 54656 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_480
timestamp 1669390400
transform 1 0 55104 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_507
timestamp 1669390400
transform 1 0 58128 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_10
timestamp 1669390400
transform 1 0 2464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_14
timestamp 1669390400
transform 1 0 2912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_19
timestamp 1669390400
transform 1 0 3472 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_25
timestamp 1669390400
transform 1 0 4144 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_33
timestamp 1669390400
transform 1 0 5040 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_40
timestamp 1669390400
transform 1 0 5824 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_44
timestamp 1669390400
transform 1 0 6272 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_49
timestamp 1669390400
transform 1 0 6832 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_65
timestamp 1669390400
transform 1 0 8624 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_96
timestamp 1669390400
transform 1 0 12096 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_100
timestamp 1669390400
transform 1 0 12544 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_104
timestamp 1669390400
transform 1 0 12992 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_116
timestamp 1669390400
transform 1 0 14336 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_118
timestamp 1669390400
transform 1 0 14560 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_123
timestamp 1669390400
transform 1 0 15120 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_129
timestamp 1669390400
transform 1 0 15792 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_137
timestamp 1669390400
transform 1 0 16688 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_139
timestamp 1669390400
transform 1 0 16912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_142
timestamp 1669390400
transform 1 0 17248 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_146
timestamp 1669390400
transform 1 0 17696 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_185
timestamp 1669390400
transform 1 0 22064 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_216
timestamp 1669390400
transform 1 0 25536 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_280
timestamp 1669390400
transform 1 0 32704 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_284
timestamp 1669390400
transform 1 0 33152 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_286
timestamp 1669390400
transform 1 0 33376 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_316
timestamp 1669390400
transform 1 0 36736 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_326
timestamp 1669390400
transform 1 0 37856 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_330
timestamp 1669390400
transform 1 0 38304 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_334
timestamp 1669390400
transform 1 0 38752 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_336
timestamp 1669390400
transform 1 0 38976 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_366
timestamp 1669390400
transform 1 0 42336 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_370
timestamp 1669390400
transform 1 0 42784 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_386
timestamp 1669390400
transform 1 0 44576 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_395
timestamp 1669390400
transform 1 0 45584 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_403
timestamp 1669390400
transform 1 0 46480 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_411
timestamp 1669390400
transform 1 0 47376 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_444
timestamp 1669390400
transform 1 0 51072 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_448
timestamp 1669390400
transform 1 0 51520 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_495
timestamp 1669390400
transform 1 0 56784 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_503
timestamp 1669390400
transform 1 0 57680 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_507
timestamp 1669390400
transform 1 0 58128 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_17
timestamp 1669390400
transform 1 0 3248 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_25
timestamp 1669390400
transform 1 0 4144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_29
timestamp 1669390400
transform 1 0 4592 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_31
timestamp 1669390400
transform 1 0 4816 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_34
timestamp 1669390400
transform 1 0 5152 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_50
timestamp 1669390400
transform 1 0 6944 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_56
timestamp 1669390400
transform 1 0 7616 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_64
timestamp 1669390400
transform 1 0 8512 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_68
timestamp 1669390400
transform 1 0 8960 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_103
timestamp 1669390400
transform 1 0 12880 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_107
timestamp 1669390400
transform 1 0 13328 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_111
timestamp 1669390400
transform 1 0 13776 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_113
timestamp 1669390400
transform 1 0 14000 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_116
timestamp 1669390400
transform 1 0 14336 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_132
timestamp 1669390400
transform 1 0 16128 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_140
timestamp 1669390400
transform 1 0 17024 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_160
timestamp 1669390400
transform 1 0 19264 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_168
timestamp 1669390400
transform 1 0 20160 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_172
timestamp 1669390400
transform 1 0 20608 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_176
timestamp 1669390400
transform 1 0 21056 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_180
timestamp 1669390400
transform 1 0 21504 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_184
timestamp 1669390400
transform 1 0 21952 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_189
timestamp 1669390400
transform 1 0 22512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_197
timestamp 1669390400
transform 1 0 23408 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_199
timestamp 1669390400
transform 1 0 23632 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_210
timestamp 1669390400
transform 1 0 24864 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_220
timestamp 1669390400
transform 1 0 25984 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_228
timestamp 1669390400
transform 1 0 26880 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_232
timestamp 1669390400
transform 1 0 27328 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_262
timestamp 1669390400
transform 1 0 30688 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_278
timestamp 1669390400
transform 1 0 32480 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_282
timestamp 1669390400
transform 1 0 32928 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_337
timestamp 1669390400
transform 1 0 39088 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_341
timestamp 1669390400
transform 1 0 39536 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_349
timestamp 1669390400
transform 1 0 40432 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_353
timestamp 1669390400
transform 1 0 40880 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_360
timestamp 1669390400
transform 1 0 41664 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_362
timestamp 1669390400
transform 1 0 41888 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_392
timestamp 1669390400
transform 1 0 45248 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_402
timestamp 1669390400
transform 1 0 46368 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_404
timestamp 1669390400
transform 1 0 46592 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_413
timestamp 1669390400
transform 1 0 47600 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1669390400
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_436
timestamp 1669390400
transform 1 0 50176 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_440
timestamp 1669390400
transform 1 0 50624 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_444
timestamp 1669390400
transform 1 0 51072 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_507
timestamp 1669390400
transform 1 0 58128 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_32
timestamp 1669390400
transform 1 0 4928 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1669390400
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_88
timestamp 1669390400
transform 1 0 11200 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_92
timestamp 1669390400
transform 1 0 11648 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_103
timestamp 1669390400
transform 1 0 12880 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_111
timestamp 1669390400
transform 1 0 13776 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_115
timestamp 1669390400
transform 1 0 14224 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_145
timestamp 1669390400
transform 1 0 17584 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_209
timestamp 1669390400
transform 1 0 24752 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_217
timestamp 1669390400
transform 1 0 25648 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_258
timestamp 1669390400
transform 1 0 30240 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_262
timestamp 1669390400
transform 1 0 30688 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_293
timestamp 1669390400
transform 1 0 34160 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_299
timestamp 1669390400
transform 1 0 34832 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_303
timestamp 1669390400
transform 1 0 35280 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_354
timestamp 1669390400
transform 1 0 40992 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_364
timestamp 1669390400
transform 1 0 42112 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_368
timestamp 1669390400
transform 1 0 42560 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_384
timestamp 1669390400
transform 1 0 44352 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_388
timestamp 1669390400
transform 1 0 44800 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_396
timestamp 1669390400
transform 1 0 45696 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_398
timestamp 1669390400
transform 1 0 45920 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_410
timestamp 1669390400
transform 1 0 47264 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_420
timestamp 1669390400
transform 1 0 48384 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_436
timestamp 1669390400
transform 1 0 50176 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_454
timestamp 1669390400
transform 1 0 52192 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_458
timestamp 1669390400
transform 1 0 52640 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_495
timestamp 1669390400
transform 1 0 56784 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_503
timestamp 1669390400
transform 1 0 57680 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_507
timestamp 1669390400
transform 1 0 58128 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_39
timestamp 1669390400
transform 1 0 5712 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_76
timestamp 1669390400
transform 1 0 9856 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_78
timestamp 1669390400
transform 1 0 10080 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_83
timestamp 1669390400
transform 1 0 10640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_87
timestamp 1669390400
transform 1 0 11088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_90
timestamp 1669390400
transform 1 0 11424 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_94
timestamp 1669390400
transform 1 0 11872 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_97
timestamp 1669390400
transform 1 0 12208 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_128
timestamp 1669390400
transform 1 0 15680 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_134
timestamp 1669390400
transform 1 0 16352 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_138
timestamp 1669390400
transform 1 0 16800 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_195
timestamp 1669390400
transform 1 0 23184 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_199
timestamp 1669390400
transform 1 0 23632 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_207
timestamp 1669390400
transform 1 0 24528 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_211
timestamp 1669390400
transform 1 0 24976 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_225
timestamp 1669390400
transform 1 0 26544 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_277
timestamp 1669390400
transform 1 0 32368 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_281
timestamp 1669390400
transform 1 0 32816 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_316
timestamp 1669390400
transform 1 0 36736 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_324
timestamp 1669390400
transform 1 0 37632 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_408
timestamp 1669390400
transform 1 0 47040 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_412
timestamp 1669390400
transform 1 0 47488 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_416
timestamp 1669390400
transform 1 0 47936 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_418
timestamp 1669390400
transform 1 0 48160 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_442
timestamp 1669390400
transform 1 0 50848 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_452
timestamp 1669390400
transform 1 0 51968 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_462
timestamp 1669390400
transform 1 0 53088 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_494
timestamp 1669390400
transform 1 0 56672 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_507
timestamp 1669390400
transform 1 0 58128 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_18
timestamp 1669390400
transform 1 0 3360 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_26
timestamp 1669390400
transform 1 0 4256 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_32
timestamp 1669390400
transform 1 0 4928 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_41
timestamp 1669390400
transform 1 0 5936 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_57
timestamp 1669390400
transform 1 0 7728 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_65
timestamp 1669390400
transform 1 0 8624 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_69
timestamp 1669390400
transform 1 0 9072 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_99
timestamp 1669390400
transform 1 0 12432 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_138
timestamp 1669390400
transform 1 0 16800 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_142
timestamp 1669390400
transform 1 0 17248 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_150
timestamp 1669390400
transform 1 0 18144 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_154
timestamp 1669390400
transform 1 0 18592 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_160
timestamp 1669390400
transform 1 0 19264 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_195
timestamp 1669390400
transform 1 0 23184 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_199
timestamp 1669390400
transform 1 0 23632 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_229
timestamp 1669390400
transform 1 0 26992 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_235
timestamp 1669390400
transform 1 0 27664 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_239
timestamp 1669390400
transform 1 0 28112 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_245
timestamp 1669390400
transform 1 0 28784 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_261
timestamp 1669390400
transform 1 0 30576 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_265
timestamp 1669390400
transform 1 0 31024 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_278
timestamp 1669390400
transform 1 0 32480 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_284
timestamp 1669390400
transform 1 0 33152 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_292
timestamp 1669390400
transform 1 0 34048 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_303
timestamp 1669390400
transform 1 0 35280 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_351
timestamp 1669390400
transform 1 0 40656 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_357
timestamp 1669390400
transform 1 0 41328 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_359
timestamp 1669390400
transform 1 0 41552 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_403
timestamp 1669390400
transform 1 0 46480 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_411
timestamp 1669390400
transform 1 0 47376 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_415
timestamp 1669390400
transform 1 0 47824 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_422
timestamp 1669390400
transform 1 0 48608 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_438
timestamp 1669390400
transform 1 0 50400 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_442
timestamp 1669390400
transform 1 0 50848 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_450
timestamp 1669390400
transform 1 0 51744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_495
timestamp 1669390400
transform 1 0 56784 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_503
timestamp 1669390400
transform 1 0 57680 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_507
timestamp 1669390400
transform 1 0 58128 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_34
timestamp 1669390400
transform 1 0 5152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_42
timestamp 1669390400
transform 1 0 6048 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_46
timestamp 1669390400
transform 1 0 6496 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_48
timestamp 1669390400
transform 1 0 6720 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_55
timestamp 1669390400
transform 1 0 7504 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_89
timestamp 1669390400
transform 1 0 11312 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_140
timestamp 1669390400
transform 1 0 17024 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_149
timestamp 1669390400
transform 1 0 18032 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_153
timestamp 1669390400
transform 1 0 18480 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_184
timestamp 1669390400
transform 1 0 21952 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_188
timestamp 1669390400
transform 1 0 22400 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_204
timestamp 1669390400
transform 1 0 24192 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_220
timestamp 1669390400
transform 1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_228
timestamp 1669390400
transform 1 0 26880 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_230
timestamp 1669390400
transform 1 0 27104 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_260
timestamp 1669390400
transform 1 0 30464 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_276
timestamp 1669390400
transform 1 0 32256 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_302
timestamp 1669390400
transform 1 0 35168 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_339
timestamp 1669390400
transform 1 0 39312 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_345
timestamp 1669390400
transform 1 0 39984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_353
timestamp 1669390400
transform 1 0 40880 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_391
timestamp 1669390400
transform 1 0 45136 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_399
timestamp 1669390400
transform 1 0 46032 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_415
timestamp 1669390400
transform 1 0 47824 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_435
timestamp 1669390400
transform 1 0 50064 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_439
timestamp 1669390400
transform 1 0 50512 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_453
timestamp 1669390400
transform 1 0 52080 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_484
timestamp 1669390400
transform 1 0 55552 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_488
timestamp 1669390400
transform 1 0 56000 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_507
timestamp 1669390400
transform 1 0 58128 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_41
timestamp 1669390400
transform 1 0 5936 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_50
timestamp 1669390400
transform 1 0 6944 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_54
timestamp 1669390400
transform 1 0 7392 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_56
timestamp 1669390400
transform 1 0 7616 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_86
timestamp 1669390400
transform 1 0 10976 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_90
timestamp 1669390400
transform 1 0 11424 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_113
timestamp 1669390400
transform 1 0 14000 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_121
timestamp 1669390400
transform 1 0 14896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_125
timestamp 1669390400
transform 1 0 15344 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_156
timestamp 1669390400
transform 1 0 18816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_164
timestamp 1669390400
transform 1 0 19712 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_183
timestamp 1669390400
transform 1 0 21840 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_214
timestamp 1669390400
transform 1 0 25312 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_218
timestamp 1669390400
transform 1 0 25760 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_234
timestamp 1669390400
transform 1 0 27552 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_238
timestamp 1669390400
transform 1 0 28000 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_266
timestamp 1669390400
transform 1 0 31136 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_296
timestamp 1669390400
transform 1 0 34496 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_300
timestamp 1669390400
transform 1 0 34944 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_316
timestamp 1669390400
transform 1 0 36736 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_326
timestamp 1669390400
transform 1 0 37856 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_332
timestamp 1669390400
transform 1 0 38528 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_340
timestamp 1669390400
transform 1 0 39424 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_373
timestamp 1669390400
transform 1 0 43120 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_377
timestamp 1669390400
transform 1 0 43568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_381
timestamp 1669390400
transform 1 0 44016 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_406
timestamp 1669390400
transform 1 0 46816 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_414
timestamp 1669390400
transform 1 0 47712 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_418
timestamp 1669390400
transform 1 0 48160 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_425
timestamp 1669390400
transform 1 0 48944 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_436
timestamp 1669390400
transform 1 0 50176 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_440
timestamp 1669390400
transform 1 0 50624 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_458
timestamp 1669390400
transform 1 0 52640 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_495
timestamp 1669390400
transform 1 0 56784 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_503
timestamp 1669390400
transform 1 0 57680 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_507
timestamp 1669390400
transform 1 0 58128 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_10
timestamp 1669390400
transform 1 0 2464 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_14
timestamp 1669390400
transform 1 0 2912 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_16
timestamp 1669390400
transform 1 0 3136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_46
timestamp 1669390400
transform 1 0 6496 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_50
timestamp 1669390400
transform 1 0 6944 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_60
timestamp 1669390400
transform 1 0 8064 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_80
timestamp 1669390400
transform 1 0 10304 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_88
timestamp 1669390400
transform 1 0 11200 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_93
timestamp 1669390400
transform 1 0 11760 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_125
timestamp 1669390400
transform 1 0 15344 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_174
timestamp 1669390400
transform 1 0 20832 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_178
timestamp 1669390400
transform 1 0 21280 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_231
timestamp 1669390400
transform 1 0 27216 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_239
timestamp 1669390400
transform 1 0 28112 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_270
timestamp 1669390400
transform 1 0 31584 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_274
timestamp 1669390400
transform 1 0 32032 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_280
timestamp 1669390400
transform 1 0 32704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_291
timestamp 1669390400
transform 1 0 33936 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_299
timestamp 1669390400
transform 1 0 34832 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_303
timestamp 1669390400
transform 1 0 35280 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_368
timestamp 1669390400
transform 1 0 42560 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_372
timestamp 1669390400
transform 1 0 43008 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_374
timestamp 1669390400
transform 1 0 43232 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_404
timestamp 1669390400
transform 1 0 46592 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_408
timestamp 1669390400
transform 1 0 47040 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_414
timestamp 1669390400
transform 1 0 47712 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_424
timestamp 1669390400
transform 1 0 48832 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_439
timestamp 1669390400
transform 1 0 50512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_443
timestamp 1669390400
transform 1 0 50960 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_449
timestamp 1669390400
transform 1 0 51632 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_457
timestamp 1669390400
transform 1 0 52528 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_461
timestamp 1669390400
transform 1 0 52976 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_464
timestamp 1669390400
transform 1 0 53312 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_472
timestamp 1669390400
transform 1 0 54208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_476
timestamp 1669390400
transform 1 0 54656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_491
timestamp 1669390400
transform 1 0 56336 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_495
timestamp 1669390400
transform 1 0 56784 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_507
timestamp 1669390400
transform 1 0 58128 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_41
timestamp 1669390400
transform 1 0 5936 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_51
timestamp 1669390400
transform 1 0 7056 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_59
timestamp 1669390400
transform 1 0 7952 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_66
timestamp 1669390400
transform 1 0 8736 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_70
timestamp 1669390400
transform 1 0 9184 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_74
timestamp 1669390400
transform 1 0 9632 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_111
timestamp 1669390400
transform 1 0 13776 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_115
timestamp 1669390400
transform 1 0 14224 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_127
timestamp 1669390400
transform 1 0 15568 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_143
timestamp 1669390400
transform 1 0 17360 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_147
timestamp 1669390400
transform 1 0 17808 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_153
timestamp 1669390400
transform 1 0 18480 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_169
timestamp 1669390400
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_173
timestamp 1669390400
transform 1 0 20720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_187
timestamp 1669390400
transform 1 0 22288 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_191
timestamp 1669390400
transform 1 0 22736 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_193
timestamp 1669390400
transform 1 0 22960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_198
timestamp 1669390400
transform 1 0 23520 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_206
timestamp 1669390400
transform 1 0 24416 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_237
timestamp 1669390400
transform 1 0 27888 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_241
timestamp 1669390400
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_245
timestamp 1669390400
transform 1 0 28784 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_266
timestamp 1669390400
transform 1 0 31136 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_274
timestamp 1669390400
transform 1 0 32032 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_304
timestamp 1669390400
transform 1 0 35392 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_312
timestamp 1669390400
transform 1 0 36288 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_316
timestamp 1669390400
transform 1 0 36736 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_354
timestamp 1669390400
transform 1 0 40992 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_368
timestamp 1669390400
transform 1 0 42560 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_384
timestamp 1669390400
transform 1 0 44352 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_388
timestamp 1669390400
transform 1 0 44800 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_400
timestamp 1669390400
transform 1 0 46144 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_430
timestamp 1669390400
transform 1 0 49504 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_442
timestamp 1669390400
transform 1 0 50848 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_452
timestamp 1669390400
transform 1 0 51968 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_458
timestamp 1669390400
transform 1 0 52640 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_496
timestamp 1669390400
transform 1 0 56896 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_504
timestamp 1669390400
transform 1 0 57792 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_508
timestamp 1669390400
transform 1 0 58240 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_34
timestamp 1669390400
transform 1 0 5152 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_38
timestamp 1669390400
transform 1 0 5600 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_40
timestamp 1669390400
transform 1 0 5824 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_47
timestamp 1669390400
transform 1 0 6608 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_63
timestamp 1669390400
transform 1 0 8400 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_89
timestamp 1669390400
transform 1 0 11312 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_97
timestamp 1669390400
transform 1 0 12208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_101
timestamp 1669390400
transform 1 0 12656 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_131
timestamp 1669390400
transform 1 0 16016 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_135
timestamp 1669390400
transform 1 0 16464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_139
timestamp 1669390400
transform 1 0 16912 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_160
timestamp 1669390400
transform 1 0 19264 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_168
timestamp 1669390400
transform 1 0 20160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_183
timestamp 1669390400
transform 1 0 21840 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_187
timestamp 1669390400
transform 1 0 22288 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_192
timestamp 1669390400
transform 1 0 22848 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_266
timestamp 1669390400
transform 1 0 31136 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_278
timestamp 1669390400
transform 1 0 32480 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_282
timestamp 1669390400
transform 1 0 32928 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_290
timestamp 1669390400
transform 1 0 33824 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_292
timestamp 1669390400
transform 1 0 34048 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_297
timestamp 1669390400
transform 1 0 34608 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_301
timestamp 1669390400
transform 1 0 35056 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_331
timestamp 1669390400
transform 1 0 38416 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_347
timestamp 1669390400
transform 1 0 40208 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_362
timestamp 1669390400
transform 1 0 41888 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_370
timestamp 1669390400
transform 1 0 42784 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_403
timestamp 1669390400
transform 1 0 46480 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_407
timestamp 1669390400
transform 1 0 46928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_415
timestamp 1669390400
transform 1 0 47824 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_419
timestamp 1669390400
transform 1 0 48272 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1669390400
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_479
timestamp 1669390400
transform 1 0 54992 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_495
timestamp 1669390400
transform 1 0 56784 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_507
timestamp 1669390400
transform 1 0 58128 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_39
timestamp 1669390400
transform 1 0 5712 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_48
timestamp 1669390400
transform 1 0 6720 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_50
timestamp 1669390400
transform 1 0 6944 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_57
timestamp 1669390400
transform 1 0 7728 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_73
timestamp 1669390400
transform 1 0 9520 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_75
timestamp 1669390400
transform 1 0 9744 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_114
timestamp 1669390400
transform 1 0 14112 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_122
timestamp 1669390400
transform 1 0 15008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_130
timestamp 1669390400
transform 1 0 15904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_134
timestamp 1669390400
transform 1 0 16352 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_164
timestamp 1669390400
transform 1 0 19712 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_168
timestamp 1669390400
transform 1 0 20160 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_183
timestamp 1669390400
transform 1 0 21840 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_199
timestamp 1669390400
transform 1 0 23632 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_207
timestamp 1669390400
transform 1 0 24528 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_209
timestamp 1669390400
transform 1 0 24752 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_214
timestamp 1669390400
transform 1 0 25312 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_226
timestamp 1669390400
transform 1 0 26656 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_234
timestamp 1669390400
transform 1 0 27552 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_238
timestamp 1669390400
transform 1 0 28000 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_241
timestamp 1669390400
transform 1 0 28336 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_304
timestamp 1669390400
transform 1 0 35392 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_308
timestamp 1669390400
transform 1 0 35840 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_310
timestamp 1669390400
transform 1 0 36064 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_315
timestamp 1669390400
transform 1 0 36624 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_329
timestamp 1669390400
transform 1 0 38192 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_333
timestamp 1669390400
transform 1 0 38640 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_338
timestamp 1669390400
transform 1 0 39200 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_354
timestamp 1669390400
transform 1 0 40992 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_362
timestamp 1669390400
transform 1 0 41888 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_367
timestamp 1669390400
transform 1 0 42448 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_375
timestamp 1669390400
transform 1 0 43344 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_379
timestamp 1669390400
transform 1 0 43792 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_381
timestamp 1669390400
transform 1 0 44016 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_386
timestamp 1669390400
transform 1 0 44576 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_424
timestamp 1669390400
transform 1 0 48832 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_426
timestamp 1669390400
transform 1 0 49056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_429
timestamp 1669390400
transform 1 0 49392 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_466
timestamp 1669390400
transform 1 0 53536 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_498
timestamp 1669390400
transform 1 0 57120 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_506
timestamp 1669390400
transform 1 0 58016 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_508
timestamp 1669390400
transform 1 0 58240 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_18
timestamp 1669390400
transform 1 0 3360 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_26
timestamp 1669390400
transform 1 0 4256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_30
timestamp 1669390400
transform 1 0 4704 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_32
timestamp 1669390400
transform 1 0 4928 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_39
timestamp 1669390400
transform 1 0 5712 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_76
timestamp 1669390400
transform 1 0 9856 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_84
timestamp 1669390400
transform 1 0 10752 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_88
timestamp 1669390400
transform 1 0 11200 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_94
timestamp 1669390400
transform 1 0 11872 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_102
timestamp 1669390400
transform 1 0 12768 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_104
timestamp 1669390400
transform 1 0 12992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_107
timestamp 1669390400
transform 1 0 13328 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_123
timestamp 1669390400
transform 1 0 15120 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_131
timestamp 1669390400
transform 1 0 16016 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_135
timestamp 1669390400
transform 1 0 16464 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_149
timestamp 1669390400
transform 1 0 18032 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_151
timestamp 1669390400
transform 1 0 18256 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_181
timestamp 1669390400
transform 1 0 21616 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_252
timestamp 1669390400
transform 1 0 29568 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_316
timestamp 1669390400
transform 1 0 36736 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_320
timestamp 1669390400
transform 1 0 37184 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_328
timestamp 1669390400
transform 1 0 38080 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_332
timestamp 1669390400
transform 1 0 38528 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_334
timestamp 1669390400
transform 1 0 38752 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_345
timestamp 1669390400
transform 1 0 39984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_349
timestamp 1669390400
transform 1 0 40432 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_351
timestamp 1669390400
transform 1 0 40656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_387
timestamp 1669390400
transform 1 0 44688 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_389
timestamp 1669390400
transform 1 0 44912 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_400
timestamp 1669390400
transform 1 0 46144 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_406
timestamp 1669390400
transform 1 0 46816 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_422
timestamp 1669390400
transform 1 0 48608 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_437
timestamp 1669390400
transform 1 0 50288 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_469
timestamp 1669390400
transform 1 0 53872 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_485
timestamp 1669390400
transform 1 0 55664 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_493
timestamp 1669390400
transform 1 0 56560 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_507
timestamp 1669390400
transform 1 0 58128 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_47
timestamp 1669390400
transform 1 0 6608 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_79
timestamp 1669390400
transform 1 0 10192 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_95
timestamp 1669390400
transform 1 0 11984 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_103
timestamp 1669390400
transform 1 0 12880 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_114
timestamp 1669390400
transform 1 0 14112 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_122
timestamp 1669390400
transform 1 0 15008 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_126
timestamp 1669390400
transform 1 0 15456 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_130
timestamp 1669390400
transform 1 0 15904 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_161
timestamp 1669390400
transform 1 0 19376 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_175
timestamp 1669390400
transform 1 0 20944 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_183
timestamp 1669390400
transform 1 0 21840 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_191
timestamp 1669390400
transform 1 0 22736 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_199
timestamp 1669390400
transform 1 0 23632 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_207
timestamp 1669390400
transform 1 0 24528 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_212
timestamp 1669390400
transform 1 0 25088 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_228
timestamp 1669390400
transform 1 0 26880 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_236
timestamp 1669390400
transform 1 0 27776 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_242
timestamp 1669390400
transform 1 0 28448 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_246
timestamp 1669390400
transform 1 0 28896 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_258
timestamp 1669390400
transform 1 0 30240 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_262
timestamp 1669390400
transform 1 0 30688 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_274
timestamp 1669390400
transform 1 0 32032 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_278
timestamp 1669390400
transform 1 0 32480 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_282
timestamp 1669390400
transform 1 0 32928 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_284
timestamp 1669390400
transform 1 0 33152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_287
timestamp 1669390400
transform 1 0 33488 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_289
timestamp 1669390400
transform 1 0 33712 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_294
timestamp 1669390400
transform 1 0 34272 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_310
timestamp 1669390400
transform 1 0 36064 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_373
timestamp 1669390400
transform 1 0 43120 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_379
timestamp 1669390400
transform 1 0 43792 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_383
timestamp 1669390400
transform 1 0 44240 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_387
timestamp 1669390400
transform 1 0 44688 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_423
timestamp 1669390400
transform 1 0 48720 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_435
timestamp 1669390400
transform 1 0 50064 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_451
timestamp 1669390400
transform 1 0 51856 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_459
timestamp 1669390400
transform 1 0 52752 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_495
timestamp 1669390400
transform 1 0 56784 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_503
timestamp 1669390400
transform 1 0 57680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_507
timestamp 1669390400
transform 1 0 58128 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_10
timestamp 1669390400
transform 1 0 2464 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_43
timestamp 1669390400
transform 1 0 6160 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_47
timestamp 1669390400
transform 1 0 6608 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_63
timestamp 1669390400
transform 1 0 8400 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_124
timestamp 1669390400
transform 1 0 15232 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_136
timestamp 1669390400
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_140
timestamp 1669390400
transform 1 0 17024 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_152
timestamp 1669390400
transform 1 0 18368 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_155
timestamp 1669390400
transform 1 0 18704 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_207
timestamp 1669390400
transform 1 0 24528 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_211
timestamp 1669390400
transform 1 0 24976 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_219
timestamp 1669390400
transform 1 0 25872 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_231
timestamp 1669390400
transform 1 0 27216 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_247
timestamp 1669390400
transform 1 0 29008 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_280
timestamp 1669390400
transform 1 0 32704 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_316
timestamp 1669390400
transform 1 0 36736 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_347
timestamp 1669390400
transform 1 0 40208 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_351
timestamp 1669390400
transform 1 0 40656 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_387
timestamp 1669390400
transform 1 0 44688 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_391
timestamp 1669390400
transform 1 0 45136 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_395
timestamp 1669390400
transform 1 0 45584 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_458
timestamp 1669390400
transform 1 0 52640 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_490
timestamp 1669390400
transform 1 0 56224 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_494
timestamp 1669390400
transform 1 0 56672 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_507
timestamp 1669390400
transform 1 0 58128 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_69
timestamp 1669390400
transform 1 0 9072 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_73
timestamp 1669390400
transform 1 0 9520 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_75
timestamp 1669390400
transform 1 0 9744 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_138
timestamp 1669390400
transform 1 0 16800 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_142
timestamp 1669390400
transform 1 0 17248 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_146
timestamp 1669390400
transform 1 0 17696 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_148
timestamp 1669390400
transform 1 0 17920 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_153
timestamp 1669390400
transform 1 0 18480 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_163
timestamp 1669390400
transform 1 0 19600 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_167
timestamp 1669390400
transform 1 0 20048 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_183
timestamp 1669390400
transform 1 0 21840 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_199
timestamp 1669390400
transform 1 0 23632 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_230
timestamp 1669390400
transform 1 0 27104 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_234
timestamp 1669390400
transform 1 0 27552 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_242
timestamp 1669390400
transform 1 0 28448 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_246
timestamp 1669390400
transform 1 0 28896 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_266
timestamp 1669390400
transform 1 0 31136 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_270
timestamp 1669390400
transform 1 0 31584 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_300
timestamp 1669390400
transform 1 0 34944 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_304
timestamp 1669390400
transform 1 0 35392 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_312
timestamp 1669390400
transform 1 0 36288 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_351
timestamp 1669390400
transform 1 0 40656 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_355
timestamp 1669390400
transform 1 0 41104 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_371
timestamp 1669390400
transform 1 0 42896 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_375
timestamp 1669390400
transform 1 0 43344 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_377
timestamp 1669390400
transform 1 0 43568 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_382
timestamp 1669390400
transform 1 0 44128 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_400
timestamp 1669390400
transform 1 0 46144 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_404
timestamp 1669390400
transform 1 0 46592 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_408
timestamp 1669390400
transform 1 0 47040 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_495
timestamp 1669390400
transform 1 0 56784 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_503
timestamp 1669390400
transform 1 0 57680 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_507
timestamp 1669390400
transform 1 0 58128 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_89
timestamp 1669390400
transform 1 0 11312 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_99
timestamp 1669390400
transform 1 0 12432 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_130
timestamp 1669390400
transform 1 0 15904 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_134
timestamp 1669390400
transform 1 0 16352 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_174
timestamp 1669390400
transform 1 0 20832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_178
timestamp 1669390400
transform 1 0 21280 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_182
timestamp 1669390400
transform 1 0 21728 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_219
timestamp 1669390400
transform 1 0 25872 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_250
timestamp 1669390400
transform 1 0 29344 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_254
timestamp 1669390400
transform 1 0 29792 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_270
timestamp 1669390400
transform 1 0 31584 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_278
timestamp 1669390400
transform 1 0 32480 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_282
timestamp 1669390400
transform 1 0 32928 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_291
timestamp 1669390400
transform 1 0 33936 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_299
timestamp 1669390400
transform 1 0 34832 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_303
timestamp 1669390400
transform 1 0 35280 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_305
timestamp 1669390400
transform 1 0 35504 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_316
timestamp 1669390400
transform 1 0 36736 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_324
timestamp 1669390400
transform 1 0 37632 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_329
timestamp 1669390400
transform 1 0 38192 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_345
timestamp 1669390400
transform 1 0 39984 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_353
timestamp 1669390400
transform 1 0 40880 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_365
timestamp 1669390400
transform 1 0 42224 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_398
timestamp 1669390400
transform 1 0 45920 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_402
timestamp 1669390400
transform 1 0 46368 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_404
timestamp 1669390400
transform 1 0 46592 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_409
timestamp 1669390400
transform 1 0 47152 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1669390400
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_430
timestamp 1669390400
transform 1 0 49504 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_435
timestamp 1669390400
transform 1 0 50064 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_467
timestamp 1669390400
transform 1 0 53648 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_483
timestamp 1669390400
transform 1 0 55440 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_491
timestamp 1669390400
transform 1 0 56336 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_495
timestamp 1669390400
transform 1 0 56784 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_507
timestamp 1669390400
transform 1 0 58128 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_45
timestamp 1669390400
transform 1 0 6384 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_49
timestamp 1669390400
transform 1 0 6832 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_54
timestamp 1669390400
transform 1 0 7392 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_86
timestamp 1669390400
transform 1 0 10976 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_91
timestamp 1669390400
transform 1 0 11536 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_99
timestamp 1669390400
transform 1 0 12432 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_103
timestamp 1669390400
transform 1 0 12880 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_113
timestamp 1669390400
transform 1 0 14000 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_144
timestamp 1669390400
transform 1 0 17472 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_175
timestamp 1669390400
transform 1 0 20944 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_184
timestamp 1669390400
transform 1 0 21952 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_196
timestamp 1669390400
transform 1 0 23296 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_227
timestamp 1669390400
transform 1 0 26768 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_233
timestamp 1669390400
transform 1 0 27440 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_237
timestamp 1669390400
transform 1 0 27888 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_245
timestamp 1669390400
transform 1 0 28784 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_258
timestamp 1669390400
transform 1 0 30240 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_262
timestamp 1669390400
transform 1 0 30688 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_337
timestamp 1669390400
transform 1 0 39088 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_345
timestamp 1669390400
transform 1 0 39984 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_347
timestamp 1669390400
transform 1 0 40208 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_377
timestamp 1669390400
transform 1 0 43568 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_381
timestamp 1669390400
transform 1 0 44016 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_398
timestamp 1669390400
transform 1 0 45920 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_430
timestamp 1669390400
transform 1 0 49504 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_446
timestamp 1669390400
transform 1 0 51296 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_454
timestamp 1669390400
transform 1 0 52192 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_458
timestamp 1669390400
transform 1 0 52640 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_495
timestamp 1669390400
transform 1 0 56784 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_503
timestamp 1669390400
transform 1 0 57680 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_507
timestamp 1669390400
transform 1 0 58128 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_34
timestamp 1669390400
transform 1 0 5152 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_38
timestamp 1669390400
transform 1 0 5600 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_40
timestamp 1669390400
transform 1 0 5824 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_76
timestamp 1669390400
transform 1 0 9856 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_84
timestamp 1669390400
transform 1 0 10752 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_88
timestamp 1669390400
transform 1 0 11200 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_140
timestamp 1669390400
transform 1 0 17024 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_149
timestamp 1669390400
transform 1 0 18032 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_153
timestamp 1669390400
transform 1 0 18480 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_157
timestamp 1669390400
transform 1 0 18928 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_161
timestamp 1669390400
transform 1 0 19376 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_191
timestamp 1669390400
transform 1 0 22736 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_195
timestamp 1669390400
transform 1 0 23184 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_211
timestamp 1669390400
transform 1 0 24976 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_247
timestamp 1669390400
transform 1 0 29008 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_277
timestamp 1669390400
transform 1 0 32368 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_281
timestamp 1669390400
transform 1 0 32816 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_288
timestamp 1669390400
transform 1 0 33600 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_293
timestamp 1669390400
transform 1 0 34160 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_301
timestamp 1669390400
transform 1 0 35056 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_331
timestamp 1669390400
transform 1 0 38416 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_333
timestamp 1669390400
transform 1 0 38640 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_338
timestamp 1669390400
transform 1 0 39200 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_342
timestamp 1669390400
transform 1 0 39648 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_411
timestamp 1669390400
transform 1 0 47376 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_417
timestamp 1669390400
transform 1 0 48048 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1669390400
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_507
timestamp 1669390400
transform 1 0 58128 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_112
timestamp 1669390400
transform 1 0 13888 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_164
timestamp 1669390400
transform 1 0 19712 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_183
timestamp 1669390400
transform 1 0 21840 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_185
timestamp 1669390400
transform 1 0 22064 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_196
timestamp 1669390400
transform 1 0 23296 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_204
timestamp 1669390400
transform 1 0 24192 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_206
timestamp 1669390400
transform 1 0 24416 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_211
timestamp 1669390400
transform 1 0 24976 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_254
timestamp 1669390400
transform 1 0 29792 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_260
timestamp 1669390400
transform 1 0 30464 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_276
timestamp 1669390400
transform 1 0 32256 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_280
timestamp 1669390400
transform 1 0 32704 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_310
timestamp 1669390400
transform 1 0 36064 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_316
timestamp 1669390400
transform 1 0 36736 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_354
timestamp 1669390400
transform 1 0 40992 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_358
timestamp 1669390400
transform 1 0 41440 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_395
timestamp 1669390400
transform 1 0 45584 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_397
timestamp 1669390400
transform 1 0 45808 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_427
timestamp 1669390400
transform 1 0 49168 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_459
timestamp 1669390400
transform 1 0 52752 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_495
timestamp 1669390400
transform 1 0 56784 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_503
timestamp 1669390400
transform 1 0 57680 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_507
timestamp 1669390400
transform 1 0 58128 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_18
timestamp 1669390400
transform 1 0 3360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_55
timestamp 1669390400
transform 1 0 7504 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_59
timestamp 1669390400
transform 1 0 7952 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_67
timestamp 1669390400
transform 1 0 8848 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_134
timestamp 1669390400
transform 1 0 16352 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_138
timestamp 1669390400
transform 1 0 16800 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_147
timestamp 1669390400
transform 1 0 17808 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_159
timestamp 1669390400
transform 1 0 19152 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_167
timestamp 1669390400
transform 1 0 20048 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_204
timestamp 1669390400
transform 1 0 24192 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_231
timestamp 1669390400
transform 1 0 27216 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_239
timestamp 1669390400
transform 1 0 28112 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_241
timestamp 1669390400
transform 1 0 28336 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_271
timestamp 1669390400
transform 1 0 31696 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_275
timestamp 1669390400
transform 1 0 32144 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_302
timestamp 1669390400
transform 1 0 35168 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_312
timestamp 1669390400
transform 1 0 36288 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_344
timestamp 1669390400
transform 1 0 39872 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_346
timestamp 1669390400
transform 1 0 40096 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_351
timestamp 1669390400
transform 1 0 40656 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_360
timestamp 1669390400
transform 1 0 41664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_364
timestamp 1669390400
transform 1 0 42112 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_415
timestamp 1669390400
transform 1 0 47824 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_419
timestamp 1669390400
transform 1 0 48272 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_423
timestamp 1669390400
transform 1 0 48720 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1669390400
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1669390400
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_507
timestamp 1669390400
transform 1 0 58128 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_42
timestamp 1669390400
transform 1 0 6048 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_48
timestamp 1669390400
transform 1 0 6720 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_52
timestamp 1669390400
transform 1 0 7168 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_66
timestamp 1669390400
transform 1 0 8736 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_97
timestamp 1669390400
transform 1 0 12208 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_114
timestamp 1669390400
transform 1 0 14112 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_145
timestamp 1669390400
transform 1 0 17584 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_187
timestamp 1669390400
transform 1 0 22288 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_203
timestamp 1669390400
transform 1 0 24080 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_205
timestamp 1669390400
transform 1 0 24304 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_235
timestamp 1669390400
transform 1 0 27664 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_239
timestamp 1669390400
transform 1 0 28112 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_255
timestamp 1669390400
transform 1 0 29904 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_287
timestamp 1669390400
transform 1 0 33488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_295
timestamp 1669390400
transform 1 0 34384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_299
timestamp 1669390400
transform 1 0 34832 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_301
timestamp 1669390400
transform 1 0 35056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_304
timestamp 1669390400
transform 1 0 35392 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_312
timestamp 1669390400
transform 1 0 36288 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_316
timestamp 1669390400
transform 1 0 36736 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_324
timestamp 1669390400
transform 1 0 37632 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_332
timestamp 1669390400
transform 1 0 38528 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_336
timestamp 1669390400
transform 1 0 38976 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_367
timestamp 1669390400
transform 1 0 42448 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_369
timestamp 1669390400
transform 1 0 42672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_380
timestamp 1669390400
transform 1 0 43904 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_386
timestamp 1669390400
transform 1 0 44576 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_396
timestamp 1669390400
transform 1 0 45696 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_427
timestamp 1669390400
transform 1 0 49168 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1669390400
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_495
timestamp 1669390400
transform 1 0 56784 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_503
timestamp 1669390400
transform 1 0 57680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_507
timestamp 1669390400
transform 1 0 58128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_34
timestamp 1669390400
transform 1 0 5152 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_64
timestamp 1669390400
transform 1 0 8512 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_68
timestamp 1669390400
transform 1 0 8960 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1669390400
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_75
timestamp 1669390400
transform 1 0 9744 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_80
timestamp 1669390400
transform 1 0 10304 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_90
timestamp 1669390400
transform 1 0 11424 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_121
timestamp 1669390400
transform 1 0 14896 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_133
timestamp 1669390400
transform 1 0 16240 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_147
timestamp 1669390400
transform 1 0 17808 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_179
timestamp 1669390400
transform 1 0 21392 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_195
timestamp 1669390400
transform 1 0 23184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_203
timestamp 1669390400
transform 1 0 24080 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_206
timestamp 1669390400
transform 1 0 24416 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_266
timestamp 1669390400
transform 1 0 31136 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_280
timestamp 1669390400
transform 1 0 32704 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_288
timestamp 1669390400
transform 1 0 33600 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_318
timestamp 1669390400
transform 1 0 36960 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_331
timestamp 1669390400
transform 1 0 38416 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_347
timestamp 1669390400
transform 1 0 40208 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_353
timestamp 1669390400
transform 1 0 40880 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_360
timestamp 1669390400
transform 1 0 41664 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_364
timestamp 1669390400
transform 1 0 42112 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_367
timestamp 1669390400
transform 1 0 42448 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_398
timestamp 1669390400
transform 1 0 45920 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_402
timestamp 1669390400
transform 1 0 46368 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_410
timestamp 1669390400
transform 1 0 47264 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_414
timestamp 1669390400
transform 1 0 47712 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_424
timestamp 1669390400
transform 1 0 48832 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_437
timestamp 1669390400
transform 1 0 50288 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_441
timestamp 1669390400
transform 1 0 50736 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_450
timestamp 1669390400
transform 1 0 51744 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_462
timestamp 1669390400
transform 1 0 53088 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_470
timestamp 1669390400
transform 1 0 53984 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_486
timestamp 1669390400
transform 1 0 55776 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_494
timestamp 1669390400
transform 1 0 56672 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1669390400
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_507
timestamp 1669390400
transform 1 0 58128 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_45
timestamp 1669390400
transform 1 0 6384 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_99
timestamp 1669390400
transform 1 0 12432 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_103
timestamp 1669390400
transform 1 0 12880 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_124
timestamp 1669390400
transform 1 0 15232 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_135
timestamp 1669390400
transform 1 0 16464 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_167
timestamp 1669390400
transform 1 0 20048 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_175
timestamp 1669390400
transform 1 0 20944 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_195
timestamp 1669390400
transform 1 0 23184 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_203
timestamp 1669390400
transform 1 0 24080 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_205
timestamp 1669390400
transform 1 0 24304 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_235
timestamp 1669390400
transform 1 0 27664 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_239
timestamp 1669390400
transform 1 0 28112 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_255
timestamp 1669390400
transform 1 0 29904 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_257
timestamp 1669390400
transform 1 0 30128 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_262
timestamp 1669390400
transform 1 0 30688 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_270
timestamp 1669390400
transform 1 0 31584 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_272
timestamp 1669390400
transform 1 0 31808 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_302
timestamp 1669390400
transform 1 0 35168 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_308
timestamp 1669390400
transform 1 0 35840 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_351
timestamp 1669390400
transform 1 0 40656 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_382
timestamp 1669390400
transform 1 0 44128 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_388
timestamp 1669390400
transform 1 0 44800 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_437
timestamp 1669390400
transform 1 0 50288 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_445
timestamp 1669390400
transform 1 0 51184 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_449
timestamp 1669390400
transform 1 0 51632 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_451
timestamp 1669390400
transform 1 0 51856 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1669390400
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_493
timestamp 1669390400
transform 1 0 56560 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_18
timestamp 1669390400
transform 1 0 3360 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_26
timestamp 1669390400
transform 1 0 4256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_59
timestamp 1669390400
transform 1 0 7952 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_67
timestamp 1669390400
transform 1 0 8848 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_92
timestamp 1669390400
transform 1 0 11648 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_94
timestamp 1669390400
transform 1 0 11872 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_99
timestamp 1669390400
transform 1 0 12432 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_130
timestamp 1669390400
transform 1 0 15904 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_138
timestamp 1669390400
transform 1 0 16800 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_146
timestamp 1669390400
transform 1 0 17696 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_151
timestamp 1669390400
transform 1 0 18256 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_196
timestamp 1669390400
transform 1 0 23296 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_200
timestamp 1669390400
transform 1 0 23744 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_220
timestamp 1669390400
transform 1 0 25984 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_224
timestamp 1669390400
transform 1 0 26432 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_236
timestamp 1669390400
transform 1 0 27776 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_238
timestamp 1669390400
transform 1 0 28000 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_268
timestamp 1669390400
transform 1 0 31360 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_272
timestamp 1669390400
transform 1 0 31808 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_280
timestamp 1669390400
transform 1 0 32704 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_291
timestamp 1669390400
transform 1 0 33936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_345
timestamp 1669390400
transform 1 0 39984 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_347
timestamp 1669390400
transform 1 0 40208 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_352
timestamp 1669390400
transform 1 0 40768 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_365
timestamp 1669390400
transform 1 0 42224 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_369
timestamp 1669390400
transform 1 0 42672 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_377
timestamp 1669390400
transform 1 0 43568 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_389
timestamp 1669390400
transform 1 0 44912 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_405
timestamp 1669390400
transform 1 0 46704 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_409
timestamp 1669390400
transform 1 0 47152 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_417
timestamp 1669390400
transform 1 0 48048 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1669390400
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_437
timestamp 1669390400
transform 1 0 50288 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_441
timestamp 1669390400
transform 1 0 50736 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_443
timestamp 1669390400
transform 1 0 50960 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_452
timestamp 1669390400
transform 1 0 51968 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_454
timestamp 1669390400
transform 1 0 52192 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_457
timestamp 1669390400
transform 1 0 52528 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_467
timestamp 1669390400
transform 1 0 53648 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_475
timestamp 1669390400
transform 1 0 54544 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_491
timestamp 1669390400
transform 1 0 56336 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_495
timestamp 1669390400
transform 1 0 56784 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_507
timestamp 1669390400
transform 1 0 58128 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_53
timestamp 1669390400
transform 1 0 7280 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_83
timestamp 1669390400
transform 1 0 10640 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_87
timestamp 1669390400
transform 1 0 11088 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_95
timestamp 1669390400
transform 1 0 11984 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_114
timestamp 1669390400
transform 1 0 14112 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_130
timestamp 1669390400
transform 1 0 15904 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_138
timestamp 1669390400
transform 1 0 16800 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_168
timestamp 1669390400
transform 1 0 20160 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_182
timestamp 1669390400
transform 1 0 21728 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_184
timestamp 1669390400
transform 1 0 21952 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_214
timestamp 1669390400
transform 1 0 25312 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_245
timestamp 1669390400
transform 1 0 28784 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_280
timestamp 1669390400
transform 1 0 32704 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_284
timestamp 1669390400
transform 1 0 33152 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_316
timestamp 1669390400
transform 1 0 36736 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_326
timestamp 1669390400
transform 1 0 37856 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_342
timestamp 1669390400
transform 1 0 39648 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_344
timestamp 1669390400
transform 1 0 39872 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_347
timestamp 1669390400
transform 1 0 40208 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_351
timestamp 1669390400
transform 1 0 40656 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_381
timestamp 1669390400
transform 1 0 44016 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_397
timestamp 1669390400
transform 1 0 45808 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_405
timestamp 1669390400
transform 1 0 46704 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_408
timestamp 1669390400
transform 1 0 47040 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1669390400
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_470
timestamp 1669390400
transform 1 0 53984 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_502
timestamp 1669390400
transform 1 0 57568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_506
timestamp 1669390400
transform 1 0 58016 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_508
timestamp 1669390400
transform 1 0 58240 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_34
timestamp 1669390400
transform 1 0 5152 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_38
timestamp 1669390400
transform 1 0 5600 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_43
timestamp 1669390400
transform 1 0 6160 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_61
timestamp 1669390400
transform 1 0 8176 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_69
timestamp 1669390400
transform 1 0 9072 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_78
timestamp 1669390400
transform 1 0 10080 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_86
timestamp 1669390400
transform 1 0 10976 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_90
timestamp 1669390400
transform 1 0 11424 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_94
timestamp 1669390400
transform 1 0 11872 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_125
timestamp 1669390400
transform 1 0 15344 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_146
timestamp 1669390400
transform 1 0 17696 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_151
timestamp 1669390400
transform 1 0 18256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_155
timestamp 1669390400
transform 1 0 18704 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_157
timestamp 1669390400
transform 1 0 18928 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_160
timestamp 1669390400
transform 1 0 19264 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_218
timestamp 1669390400
transform 1 0 25760 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_228
timestamp 1669390400
transform 1 0 26880 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_280
timestamp 1669390400
transform 1 0 32704 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_316
timestamp 1669390400
transform 1 0 36736 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_320
timestamp 1669390400
transform 1 0 37184 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_353
timestamp 1669390400
transform 1 0 40880 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_373
timestamp 1669390400
transform 1 0 43120 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_406
timestamp 1669390400
transform 1 0 46816 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_422
timestamp 1669390400
transform 1 0 48608 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_437
timestamp 1669390400
transform 1 0 50288 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_439
timestamp 1669390400
transform 1 0 50512 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_469
timestamp 1669390400
transform 1 0 53872 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_473
timestamp 1669390400
transform 1 0 54320 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_489
timestamp 1669390400
transform 1 0 56112 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_507
timestamp 1669390400
transform 1 0 58128 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_32
timestamp 1669390400
transform 1 0 4928 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1669390400
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_40
timestamp 1669390400
transform 1 0 5824 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_56
timestamp 1669390400
transform 1 0 7616 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_60
timestamp 1669390400
transform 1 0 8064 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_90
timestamp 1669390400
transform 1 0 11424 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_96
timestamp 1669390400
transform 1 0 12096 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_100
timestamp 1669390400
transform 1 0 12544 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_104
timestamp 1669390400
transform 1 0 12992 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_113
timestamp 1669390400
transform 1 0 14000 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_174
timestamp 1669390400
transform 1 0 20832 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_190
timestamp 1669390400
transform 1 0 22624 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_202
timestamp 1669390400
transform 1 0 23968 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_208
timestamp 1669390400
transform 1 0 24640 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_224
timestamp 1669390400
transform 1 0 26432 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_226
timestamp 1669390400
transform 1 0 26656 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_231
timestamp 1669390400
transform 1 0 27216 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_254
timestamp 1669390400
transform 1 0 29792 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_260
timestamp 1669390400
transform 1 0 30464 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_297
timestamp 1669390400
transform 1 0 34608 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_299
timestamp 1669390400
transform 1 0 34832 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_310
timestamp 1669390400
transform 1 0 36064 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1669390400
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_325
timestamp 1669390400
transform 1 0 37744 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_330
timestamp 1669390400
transform 1 0 38304 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_382
timestamp 1669390400
transform 1 0 44128 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_386
timestamp 1669390400
transform 1 0 44576 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_456
timestamp 1669390400
transform 1 0 52416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1669390400
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_495
timestamp 1669390400
transform 1 0 56784 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_503
timestamp 1669390400
transform 1 0 57680 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_507
timestamp 1669390400
transform 1 0 58128 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_10
timestamp 1669390400
transform 1 0 2464 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_15
timestamp 1669390400
transform 1 0 3024 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_23
timestamp 1669390400
transform 1 0 3920 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_29
timestamp 1669390400
transform 1 0 4592 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_43
timestamp 1669390400
transform 1 0 6160 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_47
timestamp 1669390400
transform 1 0 6608 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_52
timestamp 1669390400
transform 1 0 7168 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_68
timestamp 1669390400
transform 1 0 8960 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1669390400
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_127
timestamp 1669390400
transform 1 0 15568 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_131
timestamp 1669390400
transform 1 0 16016 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1669390400
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_189
timestamp 1669390400
transform 1 0 22512 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_193
timestamp 1669390400
transform 1 0 22960 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_209
timestamp 1669390400
transform 1 0 24752 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_222
timestamp 1669390400
transform 1 0 26208 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_226
timestamp 1669390400
transform 1 0 26656 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_242
timestamp 1669390400
transform 1 0 28448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_246
timestamp 1669390400
transform 1 0 28896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_276
timestamp 1669390400
transform 1 0 32256 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_282
timestamp 1669390400
transform 1 0 32928 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_290
timestamp 1669390400
transform 1 0 33824 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_296
timestamp 1669390400
transform 1 0 34496 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_300
timestamp 1669390400
transform 1 0 34944 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_308
timestamp 1669390400
transform 1 0 35840 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_341
timestamp 1669390400
transform 1 0 39536 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_349
timestamp 1669390400
transform 1 0 40432 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_353
timestamp 1669390400
transform 1 0 40880 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_387
timestamp 1669390400
transform 1 0 44688 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_391
timestamp 1669390400
transform 1 0 45136 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_423
timestamp 1669390400
transform 1 0 48720 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1669390400
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_432
timestamp 1669390400
transform 1 0 49728 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_462
timestamp 1669390400
transform 1 0 53088 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_466
timestamp 1669390400
transform 1 0 53536 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_482
timestamp 1669390400
transform 1 0 55328 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_490
timestamp 1669390400
transform 1 0 56224 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_494
timestamp 1669390400
transform 1 0 56672 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1669390400
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_507
timestamp 1669390400
transform 1 0 58128 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_4
timestamp 1669390400
transform 1 0 1792 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1669390400
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_39
timestamp 1669390400
transform 1 0 5712 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_69
timestamp 1669390400
transform 1 0 9072 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_73
timestamp 1669390400
transform 1 0 9520 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_75
timestamp 1669390400
transform 1 0 9744 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_111
timestamp 1669390400
transform 1 0 13776 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_113
timestamp 1669390400
transform 1 0 14000 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_122
timestamp 1669390400
transform 1 0 15008 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_153
timestamp 1669390400
transform 1 0 18480 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_157
timestamp 1669390400
transform 1 0 18928 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_165
timestamp 1669390400
transform 1 0 19824 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_167
timestamp 1669390400
transform 1 0 20048 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_195
timestamp 1669390400
transform 1 0 23184 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_226
timestamp 1669390400
transform 1 0 26656 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_242
timestamp 1669390400
transform 1 0 28448 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_246
timestamp 1669390400
transform 1 0 28896 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_282
timestamp 1669390400
transform 1 0 32928 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_286
timestamp 1669390400
transform 1 0 33376 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_316
timestamp 1669390400
transform 1 0 36736 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1669390400
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_326
timestamp 1669390400
transform 1 0 37856 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_330
timestamp 1669390400
transform 1 0 38304 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_361
timestamp 1669390400
transform 1 0 41776 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_373
timestamp 1669390400
transform 1 0 43120 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_381
timestamp 1669390400
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_385
timestamp 1669390400
transform 1 0 44464 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1669390400
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_422
timestamp 1669390400
transform 1 0 48608 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_453
timestamp 1669390400
transform 1 0 52080 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_457
timestamp 1669390400
transform 1 0 52528 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_495
timestamp 1669390400
transform 1 0 56784 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_503
timestamp 1669390400
transform 1 0 57680 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_507
timestamp 1669390400
transform 1 0 58128 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_10
timestamp 1669390400
transform 1 0 2464 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_15
timestamp 1669390400
transform 1 0 3024 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_67
timestamp 1669390400
transform 1 0 8848 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_82
timestamp 1669390400
transform 1 0 10528 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_86
timestamp 1669390400
transform 1 0 10976 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_102
timestamp 1669390400
transform 1 0 12768 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_106
timestamp 1669390400
transform 1 0 13216 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_108
timestamp 1669390400
transform 1 0 13440 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_113
timestamp 1669390400
transform 1 0 14000 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_121
timestamp 1669390400
transform 1 0 14896 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_133
timestamp 1669390400
transform 1 0 16240 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1669390400
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_148
timestamp 1669390400
transform 1 0 17920 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_179
timestamp 1669390400
transform 1 0 21392 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_183
timestamp 1669390400
transform 1 0 21840 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_199
timestamp 1669390400
transform 1 0 23632 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_207
timestamp 1669390400
transform 1 0 24528 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_211
timestamp 1669390400
transform 1 0 24976 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_229
timestamp 1669390400
transform 1 0 26992 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_233
timestamp 1669390400
transform 1 0 27440 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_264
timestamp 1669390400
transform 1 0 30912 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_268
timestamp 1669390400
transform 1 0 31360 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_338
timestamp 1669390400
transform 1 0 39200 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_340
timestamp 1669390400
transform 1 0 39424 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_345
timestamp 1669390400
transform 1 0 39984 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_349
timestamp 1669390400
transform 1 0 40432 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_353
timestamp 1669390400
transform 1 0 40880 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_361
timestamp 1669390400
transform 1 0 41776 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_413
timestamp 1669390400
transform 1 0 47600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_417
timestamp 1669390400
transform 1 0 48048 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_422
timestamp 1669390400
transform 1 0 48608 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_431
timestamp 1669390400
transform 1 0 49616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_435
timestamp 1669390400
transform 1 0 50064 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_437
timestamp 1669390400
transform 1 0 50288 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_442
timestamp 1669390400
transform 1 0 50848 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_494
timestamp 1669390400
transform 1 0 56672 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1669390400
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_507
timestamp 1669390400
transform 1 0 58128 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_32
timestamp 1669390400
transform 1 0 4928 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_39
timestamp 1669390400
transform 1 0 5712 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_42
timestamp 1669390400
transform 1 0 6048 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_73
timestamp 1669390400
transform 1 0 9520 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_82
timestamp 1669390400
transform 1 0 10528 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_98
timestamp 1669390400
transform 1 0 12320 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_138
timestamp 1669390400
transform 1 0 16800 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_142
timestamp 1669390400
transform 1 0 17248 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_158
timestamp 1669390400
transform 1 0 19040 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_163
timestamp 1669390400
transform 1 0 19600 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_171
timestamp 1669390400
transform 1 0 20496 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_173
timestamp 1669390400
transform 1 0 20720 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_210
timestamp 1669390400
transform 1 0 24864 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_224
timestamp 1669390400
transform 1 0 26432 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_234
timestamp 1669390400
transform 1 0 27552 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_242
timestamp 1669390400
transform 1 0 28448 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_244
timestamp 1669390400
transform 1 0 28672 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_259
timestamp 1669390400
transform 1 0 30352 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_267
timestamp 1669390400
transform 1 0 31248 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_283
timestamp 1669390400
transform 1 0 33040 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_287
timestamp 1669390400
transform 1 0 33488 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_293
timestamp 1669390400
transform 1 0 34160 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_309
timestamp 1669390400
transform 1 0 35952 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1669390400
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_353
timestamp 1669390400
transform 1 0 40880 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_361
timestamp 1669390400
transform 1 0 41776 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_369
timestamp 1669390400
transform 1 0 42672 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_394
timestamp 1669390400
transform 1 0 45472 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_399
timestamp 1669390400
transform 1 0 46032 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_405
timestamp 1669390400
transform 1 0 46704 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_409
timestamp 1669390400
transform 1 0 47152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_428
timestamp 1669390400
transform 1 0 49280 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_436
timestamp 1669390400
transform 1 0 50176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_440
timestamp 1669390400
transform 1 0 50624 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_444
timestamp 1669390400
transform 1 0 51072 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_452
timestamp 1669390400
transform 1 0 51968 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_456
timestamp 1669390400
transform 1 0 52416 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1669390400
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_482
timestamp 1669390400
transform 1 0 55328 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_498
timestamp 1669390400
transform 1 0 57120 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_506
timestamp 1669390400
transform 1 0 58016 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_508
timestamp 1669390400
transform 1 0 58240 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_10
timestamp 1669390400
transform 1 0 2464 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_15
timestamp 1669390400
transform 1 0 3024 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_31
timestamp 1669390400
transform 1 0 4816 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_34
timestamp 1669390400
transform 1 0 5152 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_50
timestamp 1669390400
transform 1 0 6944 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_56
timestamp 1669390400
transform 1 0 7616 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_64
timestamp 1669390400
transform 1 0 8512 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_68
timestamp 1669390400
transform 1 0 8960 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1669390400
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_83
timestamp 1669390400
transform 1 0 10640 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_99
timestamp 1669390400
transform 1 0 12432 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_107
timestamp 1669390400
transform 1 0 13328 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_115
timestamp 1669390400
transform 1 0 14224 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_131
timestamp 1669390400
transform 1 0 16016 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_133
timestamp 1669390400
transform 1 0 16240 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_136
timestamp 1669390400
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_140
timestamp 1669390400
transform 1 0 17024 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_149
timestamp 1669390400
transform 1 0 18032 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_157
timestamp 1669390400
transform 1 0 18928 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_161
timestamp 1669390400
transform 1 0 19376 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_163
timestamp 1669390400
transform 1 0 19600 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_193
timestamp 1669390400
transform 1 0 22960 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_197
timestamp 1669390400
transform 1 0 23408 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_224
timestamp 1669390400
transform 1 0 26432 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_228
timestamp 1669390400
transform 1 0 26880 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_236
timestamp 1669390400
transform 1 0 27776 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_243
timestamp 1669390400
transform 1 0 28560 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_251
timestamp 1669390400
transform 1 0 29456 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_255
timestamp 1669390400
transform 1 0 29904 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_257
timestamp 1669390400
transform 1 0 30128 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_269
timestamp 1669390400
transform 1 0 31472 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_277
timestamp 1669390400
transform 1 0 32368 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_281
timestamp 1669390400
transform 1 0 32816 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_294
timestamp 1669390400
transform 1 0 34272 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_298
timestamp 1669390400
transform 1 0 34720 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_300
timestamp 1669390400
transform 1 0 34944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_330
timestamp 1669390400
transform 1 0 38304 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_334
timestamp 1669390400
transform 1 0 38752 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_368
timestamp 1669390400
transform 1 0 42560 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_376
timestamp 1669390400
transform 1 0 43456 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_406
timestamp 1669390400
transform 1 0 46816 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_410
timestamp 1669390400
transform 1 0 47264 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_458
timestamp 1669390400
transform 1 0 52640 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_489
timestamp 1669390400
transform 1 0 56112 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_493
timestamp 1669390400
transform 1 0 56560 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_507
timestamp 1669390400
transform 1 0 58128 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_4
timestamp 1669390400
transform 1 0 1792 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1669390400
transform 1 0 5152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_40
timestamp 1669390400
transform 1 0 5824 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_56
timestamp 1669390400
transform 1 0 7616 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_62
timestamp 1669390400
transform 1 0 8288 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_72
timestamp 1669390400
transform 1 0 9408 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_76
timestamp 1669390400
transform 1 0 9856 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_78
timestamp 1669390400
transform 1 0 10080 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_87
timestamp 1669390400
transform 1 0 11088 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_111
timestamp 1669390400
transform 1 0 13776 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_115
timestamp 1669390400
transform 1 0 14224 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_145
timestamp 1669390400
transform 1 0 17584 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1669390400
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_190
timestamp 1669390400
transform 1 0 22624 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_194
timestamp 1669390400
transform 1 0 23072 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_210
timestamp 1669390400
transform 1 0 24864 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_214
timestamp 1669390400
transform 1 0 25312 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_231
timestamp 1669390400
transform 1 0 27216 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_241
timestamp 1669390400
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_260
timestamp 1669390400
transform 1 0 30464 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_291
timestamp 1669390400
transform 1 0 33936 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_295
timestamp 1669390400
transform 1 0 34384 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_311
timestamp 1669390400
transform 1 0 36176 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_351
timestamp 1669390400
transform 1 0 40656 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_382
timestamp 1669390400
transform 1 0 44128 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_386
timestamp 1669390400
transform 1 0 44576 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_422
timestamp 1669390400
transform 1 0 48608 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_426
timestamp 1669390400
transform 1 0 49056 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_434
timestamp 1669390400
transform 1 0 49952 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_450
timestamp 1669390400
transform 1 0 51744 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_456
timestamp 1669390400
transform 1 0 52416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1669390400
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_467
timestamp 1669390400
transform 1 0 53648 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_473
timestamp 1669390400
transform 1 0 54320 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_505
timestamp 1669390400
transform 1 0 57904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_22
timestamp 1669390400
transform 1 0 3808 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_30
timestamp 1669390400
transform 1 0 4704 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_60
timestamp 1669390400
transform 1 0 8064 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1669390400
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_103
timestamp 1669390400
transform 1 0 12880 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_134
timestamp 1669390400
transform 1 0 16352 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_138
timestamp 1669390400
transform 1 0 16800 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_147
timestamp 1669390400
transform 1 0 17808 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_201
timestamp 1669390400
transform 1 0 23856 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_205
timestamp 1669390400
transform 1 0 24304 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1669390400
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_224
timestamp 1669390400
transform 1 0 26432 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_230
timestamp 1669390400
transform 1 0 27104 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_238
timestamp 1669390400
transform 1 0 28000 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_269
timestamp 1669390400
transform 1 0 31472 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_273
timestamp 1669390400
transform 1 0 31920 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_281
timestamp 1669390400
transform 1 0 32816 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1669390400
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_320
timestamp 1669390400
transform 1 0 37184 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_328
timestamp 1669390400
transform 1 0 38080 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_333
timestamp 1669390400
transform 1 0 38640 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_349
timestamp 1669390400
transform 1 0 40432 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_353
timestamp 1669390400
transform 1 0 40880 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_369
timestamp 1669390400
transform 1 0 42672 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_400
timestamp 1669390400
transform 1 0 46144 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_404
timestamp 1669390400
transform 1 0 46592 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_406
timestamp 1669390400
transform 1 0 46816 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_423
timestamp 1669390400
transform 1 0 48720 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1669390400
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_431
timestamp 1669390400
transform 1 0 49616 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_439
timestamp 1669390400
transform 1 0 50512 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_443
timestamp 1669390400
transform 1 0 50960 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_473
timestamp 1669390400
transform 1 0 54320 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_477
timestamp 1669390400
transform 1 0 54768 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_493
timestamp 1669390400
transform 1 0 56560 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_507
timestamp 1669390400
transform 1 0 58128 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1669390400
transform 1 0 5152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_45
timestamp 1669390400
transform 1 0 6384 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_49
timestamp 1669390400
transform 1 0 6832 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_51
timestamp 1669390400
transform 1 0 7056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_60
timestamp 1669390400
transform 1 0 8064 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_71
timestamp 1669390400
transform 1 0 9296 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_75
timestamp 1669390400
transform 1 0 9744 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_83
timestamp 1669390400
transform 1 0 10640 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_91
timestamp 1669390400
transform 1 0 11536 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_93
timestamp 1669390400
transform 1 0 11760 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_159
timestamp 1669390400
transform 1 0 19152 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_165
timestamp 1669390400
transform 1 0 19824 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_169
timestamp 1669390400
transform 1 0 20272 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_171
timestamp 1669390400
transform 1 0 20496 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1669390400
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_188
timestamp 1669390400
transform 1 0 22400 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_208
timestamp 1669390400
transform 1 0 24640 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_239
timestamp 1669390400
transform 1 0 28112 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1669390400
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_253
timestamp 1669390400
transform 1 0 29680 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_267
timestamp 1669390400
transform 1 0 31248 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_277
timestamp 1669390400
transform 1 0 32368 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_285
timestamp 1669390400
transform 1 0 33264 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1669390400
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_332
timestamp 1669390400
transform 1 0 38528 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_340
timestamp 1669390400
transform 1 0 39424 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_372
timestamp 1669390400
transform 1 0 43008 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_388
timestamp 1669390400
transform 1 0 44800 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_399
timestamp 1669390400
transform 1 0 46032 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_407
timestamp 1669390400
transform 1 0 46928 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_437
timestamp 1669390400
transform 1 0 50288 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_441
timestamp 1669390400
transform 1 0 50736 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_449
timestamp 1669390400
transform 1 0 51632 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_451
timestamp 1669390400
transform 1 0 51856 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_456
timestamp 1669390400
transform 1 0 52416 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_460
timestamp 1669390400
transform 1 0 52864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_482
timestamp 1669390400
transform 1 0 55328 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_498
timestamp 1669390400
transform 1 0 57120 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_506
timestamp 1669390400
transform 1 0 58016 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_508
timestamp 1669390400
transform 1 0 58240 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_34
timestamp 1669390400
transform 1 0 5152 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_50
timestamp 1669390400
transform 1 0 6944 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_60
timestamp 1669390400
transform 1 0 8064 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_68
timestamp 1669390400
transform 1 0 8960 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1669390400
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_76
timestamp 1669390400
transform 1 0 9856 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_92
timestamp 1669390400
transform 1 0 11648 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_96
timestamp 1669390400
transform 1 0 12096 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_106
timestamp 1669390400
transform 1 0 13216 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_108
timestamp 1669390400
transform 1 0 13440 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_122
timestamp 1669390400
transform 1 0 15008 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_138
timestamp 1669390400
transform 1 0 16800 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_147
timestamp 1669390400
transform 1 0 17808 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_151
timestamp 1669390400
transform 1 0 18256 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_153
timestamp 1669390400
transform 1 0 18480 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_158
timestamp 1669390400
transform 1 0 19040 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_174
timestamp 1669390400
transform 1 0 20832 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_177
timestamp 1669390400
transform 1 0 21168 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_193
timestamp 1669390400
transform 1 0 22960 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_201
timestamp 1669390400
transform 1 0 23856 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_203
timestamp 1669390400
transform 1 0 24080 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_209
timestamp 1669390400
transform 1 0 24752 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_220
timestamp 1669390400
transform 1 0 25984 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_224
timestamp 1669390400
transform 1 0 26432 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_275
timestamp 1669390400
transform 1 0 32144 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1669390400
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_316
timestamp 1669390400
transform 1 0 36736 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_320
timestamp 1669390400
transform 1 0 37184 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_324
timestamp 1669390400
transform 1 0 37632 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_360
timestamp 1669390400
transform 1 0 41664 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_389
timestamp 1669390400
transform 1 0 44912 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_405
timestamp 1669390400
transform 1 0 46704 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_413
timestamp 1669390400
transform 1 0 47600 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_415
timestamp 1669390400
transform 1 0 47824 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_420
timestamp 1669390400
transform 1 0 48384 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_422
timestamp 1669390400
transform 1 0 48608 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1669390400
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_479
timestamp 1669390400
transform 1 0 54992 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_495
timestamp 1669390400
transform 1 0 56784 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_507
timestamp 1669390400
transform 1 0 58128 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1669390400
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_45
timestamp 1669390400
transform 1 0 6384 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_49
timestamp 1669390400
transform 1 0 6832 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_51
timestamp 1669390400
transform 1 0 7056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_60
timestamp 1669390400
transform 1 0 8064 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_68
timestamp 1669390400
transform 1 0 8960 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_84
timestamp 1669390400
transform 1 0 10752 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_92
timestamp 1669390400
transform 1 0 11648 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_96
timestamp 1669390400
transform 1 0 12096 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_112
timestamp 1669390400
transform 1 0 13888 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_114
timestamp 1669390400
transform 1 0 14112 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_144
timestamp 1669390400
transform 1 0 17472 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_175
timestamp 1669390400
transform 1 0 20944 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_190
timestamp 1669390400
transform 1 0 22624 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_221
timestamp 1669390400
transform 1 0 26096 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_231
timestamp 1669390400
transform 1 0 27216 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_235
timestamp 1669390400
transform 1 0 27664 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_238
timestamp 1669390400
transform 1 0 28000 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_246
timestamp 1669390400
transform 1 0 28896 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_254
timestamp 1669390400
transform 1 0 29792 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_268
timestamp 1669390400
transform 1 0 31360 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_284
timestamp 1669390400
transform 1 0 33152 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_292
timestamp 1669390400
transform 1 0 34048 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_300
timestamp 1669390400
transform 1 0 34944 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_305
timestamp 1669390400
transform 1 0 35504 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_309
timestamp 1669390400
transform 1 0 35952 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_311
timestamp 1669390400
transform 1 0 36176 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_314
timestamp 1669390400
transform 1 0 36512 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1669390400
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_351
timestamp 1669390400
transform 1 0 40656 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_382
timestamp 1669390400
transform 1 0 44128 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_399
timestamp 1669390400
transform 1 0 46032 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_407
timestamp 1669390400
transform 1 0 46928 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_411
timestamp 1669390400
transform 1 0 47376 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_419
timestamp 1669390400
transform 1 0 48272 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_427
timestamp 1669390400
transform 1 0 49168 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_458
timestamp 1669390400
transform 1 0 52640 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1669390400
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_494
timestamp 1669390400
transform 1 0 56672 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_498
timestamp 1669390400
transform 1 0 57120 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_506
timestamp 1669390400
transform 1 0 58016 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_508
timestamp 1669390400
transform 1 0 58240 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_18
timestamp 1669390400
transform 1 0 3360 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_22
timestamp 1669390400
transform 1 0 3808 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_53
timestamp 1669390400
transform 1 0 7280 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_61
timestamp 1669390400
transform 1 0 8176 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1669390400
transform 1 0 9184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_80
timestamp 1669390400
transform 1 0 10304 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_88
timestamp 1669390400
transform 1 0 11200 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_96
timestamp 1669390400
transform 1 0 12096 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_104
timestamp 1669390400
transform 1 0 12992 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_114
timestamp 1669390400
transform 1 0 14112 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_130
timestamp 1669390400
transform 1 0 15904 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_132
timestamp 1669390400
transform 1 0 16128 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1669390400
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_160
timestamp 1669390400
transform 1 0 19264 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_164
timestamp 1669390400
transform 1 0 19712 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_194
timestamp 1669390400
transform 1 0 23072 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_198
timestamp 1669390400
transform 1 0 23520 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_206
timestamp 1669390400
transform 1 0 24416 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1669390400
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_222
timestamp 1669390400
transform 1 0 26208 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_226
timestamp 1669390400
transform 1 0 26656 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_228
timestamp 1669390400
transform 1 0 26880 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_231
timestamp 1669390400
transform 1 0 27216 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_262
timestamp 1669390400
transform 1 0 30688 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_266
timestamp 1669390400
transform 1 0 31136 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_282
timestamp 1669390400
transform 1 0 32928 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_302
timestamp 1669390400
transform 1 0 35168 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_362
timestamp 1669390400
transform 1 0 41888 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_366
timestamp 1669390400
transform 1 0 42336 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_378
timestamp 1669390400
transform 1 0 43680 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_409
timestamp 1669390400
transform 1 0 47152 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_417
timestamp 1669390400
transform 1 0 48048 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_436
timestamp 1669390400
transform 1 0 50176 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_440
timestamp 1669390400
transform 1 0 50624 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_442
timestamp 1669390400
transform 1 0 50848 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_472
timestamp 1669390400
transform 1 0 54208 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_476
timestamp 1669390400
transform 1 0 54656 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_491
timestamp 1669390400
transform 1 0 56336 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_495
timestamp 1669390400
transform 1 0 56784 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_507
timestamp 1669390400
transform 1 0 58128 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_4
timestamp 1669390400
transform 1 0 1792 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1669390400
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_74
timestamp 1669390400
transform 1 0 9632 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1669390400
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_138
timestamp 1669390400
transform 1 0 16800 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_142
timestamp 1669390400
transform 1 0 17248 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_174
timestamp 1669390400
transform 1 0 20832 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1669390400
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_184
timestamp 1669390400
transform 1 0 21952 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_200
timestamp 1669390400
transform 1 0 23744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_233
timestamp 1669390400
transform 1 0 27440 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_237
timestamp 1669390400
transform 1 0 27888 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_245
timestamp 1669390400
transform 1 0 28784 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1669390400
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_282
timestamp 1669390400
transform 1 0 32928 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_302
timestamp 1669390400
transform 1 0 35168 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_326
timestamp 1669390400
transform 1 0 37856 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_334
timestamp 1669390400
transform 1 0 38752 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_338
timestamp 1669390400
transform 1 0 39200 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_342
timestamp 1669390400
transform 1 0 39648 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_373
timestamp 1669390400
transform 1 0 43120 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_424
timestamp 1669390400
transform 1 0 48832 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_427
timestamp 1669390400
transform 1 0 49168 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_439
timestamp 1669390400
transform 1 0 50512 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_455
timestamp 1669390400
transform 1 0 52304 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_459
timestamp 1669390400
transform 1 0 52752 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_466
timestamp 1669390400
transform 1 0 53536 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_470
timestamp 1669390400
transform 1 0 53984 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_474
timestamp 1669390400
transform 1 0 54432 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_506
timestamp 1669390400
transform 1 0 58016 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_508
timestamp 1669390400
transform 1 0 58240 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_18
timestamp 1669390400
transform 1 0 3360 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1669390400
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_76
timestamp 1669390400
transform 1 0 9856 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_92
timestamp 1669390400
transform 1 0 11648 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_100
timestamp 1669390400
transform 1 0 12544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_104
timestamp 1669390400
transform 1 0 12992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_107
timestamp 1669390400
transform 1 0 13328 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_139
timestamp 1669390400
transform 1 0 16912 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_181
timestamp 1669390400
transform 1 0 21616 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_185
timestamp 1669390400
transform 1 0 22064 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_201
timestamp 1669390400
transform 1 0 23856 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_209
timestamp 1669390400
transform 1 0 24752 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_219
timestamp 1669390400
transform 1 0 25872 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_223
timestamp 1669390400
transform 1 0 26320 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_255
timestamp 1669390400
transform 1 0 29904 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_271
timestamp 1669390400
transform 1 0 31696 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1669390400
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_319
timestamp 1669390400
transform 1 0 37072 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_323
timestamp 1669390400
transform 1 0 37520 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_362
timestamp 1669390400
transform 1 0 41888 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_394
timestamp 1669390400
transform 1 0 45472 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1669390400
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_458
timestamp 1669390400
transform 1 0 52640 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_462
timestamp 1669390400
transform 1 0 53088 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_494
timestamp 1669390400
transform 1 0 56672 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1669390400
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_507
timestamp 1669390400
transform 1 0 58128 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1669390400
transform 1 0 5152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_53
timestamp 1669390400
transform 1 0 7280 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_67
timestamp 1669390400
transform 1 0 8848 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_71
timestamp 1669390400
transform 1 0 9296 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_103
timestamp 1669390400
transform 1 0 12880 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_140
timestamp 1669390400
transform 1 0 17024 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_156
timestamp 1669390400
transform 1 0 18816 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_160
timestamp 1669390400
transform 1 0 19264 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_165
timestamp 1669390400
transform 1 0 19824 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_173
timestamp 1669390400
transform 1 0 20720 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1669390400
transform 1 0 28560 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1669390400
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1669390400
transform 1 0 36512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1669390400
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_385
timestamp 1669390400
transform 1 0 44464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1669390400
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_456
timestamp 1669390400
transform 1 0 52416 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_460
timestamp 1669390400
transform 1 0 52864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_495
timestamp 1669390400
transform 1 0 56784 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_503
timestamp 1669390400
transform 1 0 57680 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_507
timestamp 1669390400
transform 1 0 58128 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1669390400
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1669390400
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1669390400
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1669390400
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1669390400
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1669390400
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1669390400
transform 1 0 40544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_421
timestamp 1669390400
transform 1 0 48496 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1669390400
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_492
timestamp 1669390400
transform 1 0 56448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1669390400
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_507
timestamp 1669390400
transform 1 0 58128 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1669390400
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1669390400
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1669390400
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1669390400
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1669390400
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1669390400
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1669390400
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_385
timestamp 1669390400
transform 1 0 44464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_456
timestamp 1669390400
transform 1 0 52416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1669390400
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_495
timestamp 1669390400
transform 1 0 56784 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_503
timestamp 1669390400
transform 1 0 57680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_507
timestamp 1669390400
transform 1 0 58128 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1669390400
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1669390400
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1669390400
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1669390400
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1669390400
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1669390400
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1669390400
transform 1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_421
timestamp 1669390400
transform 1 0 48496 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1669390400
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_492
timestamp 1669390400
transform 1 0 56448 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1669390400
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_507
timestamp 1669390400
transform 1 0 58128 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1669390400
transform 1 0 5152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1669390400
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1669390400
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_172
timestamp 1669390400
transform 1 0 20608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1669390400
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_243
timestamp 1669390400
transform 1 0 28560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1669390400
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1669390400
transform 1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1669390400
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_385
timestamp 1669390400
transform 1 0 44464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1669390400
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_456
timestamp 1669390400
transform 1 0 52416 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1669390400
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_495
timestamp 1669390400
transform 1 0 56784 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_503
timestamp 1669390400
transform 1 0 57680 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_507
timestamp 1669390400
transform 1 0 58128 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_18
timestamp 1669390400
transform 1 0 3360 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_26
timestamp 1669390400
transform 1 0 4256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_30
timestamp 1669390400
transform 1 0 4704 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_34
timestamp 1669390400
transform 1 0 5152 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_37
timestamp 1669390400
transform 1 0 5488 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_52
timestamp 1669390400
transform 1 0 7168 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_68
timestamp 1669390400
transform 1 0 8960 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_72
timestamp 1669390400
transform 1 0 9408 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_104
timestamp 1669390400
transform 1 0 12992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_107
timestamp 1669390400
transform 1 0 13328 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_139
timestamp 1669390400
transform 1 0 16912 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_142
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_174
timestamp 1669390400
transform 1 0 20832 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_177
timestamp 1669390400
transform 1 0 21168 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_209
timestamp 1669390400
transform 1 0 24752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_228
timestamp 1669390400
transform 1 0 26880 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_243
timestamp 1669390400
transform 1 0 28560 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_247
timestamp 1669390400
transform 1 0 29008 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_279
timestamp 1669390400
transform 1 0 32592 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_282
timestamp 1669390400
transform 1 0 32928 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_314
timestamp 1669390400
transform 1 0 36512 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_317
timestamp 1669390400
transform 1 0 36848 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_349
timestamp 1669390400
transform 1 0 40432 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_352
timestamp 1669390400
transform 1 0 40768 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_384
timestamp 1669390400
transform 1 0 44352 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_387
timestamp 1669390400
transform 1 0 44688 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_419
timestamp 1669390400
transform 1 0 48272 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_422
timestamp 1669390400
transform 1 0 48608 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_426
timestamp 1669390400
transform 1 0 49056 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_441
timestamp 1669390400
transform 1 0 50736 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_449
timestamp 1669390400
transform 1 0 51632 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_453
timestamp 1669390400
transform 1 0 52080 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_457
timestamp 1669390400
transform 1 0 52528 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_489
timestamp 1669390400
transform 1 0 56112 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_492
timestamp 1669390400
transform 1 0 56448 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_508
timestamp 1669390400
transform 1 0 58240 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 5264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 13104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 20944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 28784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 36624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 44464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 52304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0475_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 52976 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0476_
timestamp 1669390400
transform 1 0 52976 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0477_
timestamp 1669390400
transform -1 0 54432 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0478_
timestamp 1669390400
transform 1 0 53312 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0479_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 54320 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0480_
timestamp 1669390400
transform 1 0 45472 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0481_
timestamp 1669390400
transform 1 0 45024 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0482_
timestamp 1669390400
transform 1 0 45472 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0483_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 46816 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0484_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 54096 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0485_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53312 0 1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0486_
timestamp 1669390400
transform 1 0 53312 0 1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0487_
timestamp 1669390400
transform 1 0 47264 0 1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0488_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 43680 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0489_
timestamp 1669390400
transform 1 0 37408 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0490_
timestamp 1669390400
transform 1 0 41440 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0491_
timestamp 1669390400
transform 1 0 42000 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0492_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 41440 0 -1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0493_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 48720 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0494_
timestamp 1669390400
transform 1 0 47376 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0495_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 38416 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0496_
timestamp 1669390400
transform 1 0 38192 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0497_
timestamp 1669390400
transform 1 0 33488 0 -1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0498_
timestamp 1669390400
transform 1 0 30800 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0499_
timestamp 1669390400
transform 1 0 29456 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0500_
timestamp 1669390400
transform 1 0 31360 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0501_
timestamp 1669390400
transform -1 0 35280 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0502_
timestamp 1669390400
transform 1 0 31248 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0503_
timestamp 1669390400
transform 1 0 37184 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0504_
timestamp 1669390400
transform 1 0 39648 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0505_
timestamp 1669390400
transform 1 0 14448 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0506_
timestamp 1669390400
transform -1 0 16576 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0507_
timestamp 1669390400
transform 1 0 19824 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0508_
timestamp 1669390400
transform 1 0 19936 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0509_
timestamp 1669390400
transform 1 0 25536 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0510_
timestamp 1669390400
transform -1 0 27216 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0511_
timestamp 1669390400
transform 1 0 20608 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0512_
timestamp 1669390400
transform -1 0 15904 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0513_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 8736 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0514_
timestamp 1669390400
transform 1 0 6832 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0515_
timestamp 1669390400
transform 1 0 43792 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0516_
timestamp 1669390400
transform 1 0 42784 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0517_
timestamp 1669390400
transform 1 0 34944 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0518_
timestamp 1669390400
transform 1 0 31584 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0519_
timestamp 1669390400
transform 1 0 35616 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0520_
timestamp 1669390400
transform 1 0 36064 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0521_
timestamp 1669390400
transform 1 0 37184 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0522_
timestamp 1669390400
transform 1 0 42784 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0523_
timestamp 1669390400
transform 1 0 50512 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0524_
timestamp 1669390400
transform 1 0 53312 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0525_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 18704 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0526_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22848 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0527_
timestamp 1669390400
transform 1 0 27664 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0528_
timestamp 1669390400
transform 1 0 31920 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0529_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 28784 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0530_
timestamp 1669390400
transform 1 0 21616 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0531_
timestamp 1669390400
transform 1 0 23744 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0532_
timestamp 1669390400
transform 1 0 23184 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0533_
timestamp 1669390400
transform -1 0 24528 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0534_
timestamp 1669390400
transform -1 0 21056 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0535_
timestamp 1669390400
transform 1 0 4816 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0536_
timestamp 1669390400
transform 1 0 9632 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0537_
timestamp 1669390400
transform 1 0 15344 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0538_
timestamp 1669390400
transform 1 0 15120 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0539_
timestamp 1669390400
transform -1 0 15008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0540_
timestamp 1669390400
transform 1 0 7392 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0541_
timestamp 1669390400
transform 1 0 9632 0 -1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0542_
timestamp 1669390400
transform -1 0 10528 0 1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0543_
timestamp 1669390400
transform 1 0 8176 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0544_
timestamp 1669390400
transform 1 0 21504 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0545_
timestamp 1669390400
transform 1 0 21504 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0546_
timestamp 1669390400
transform -1 0 22400 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0547_
timestamp 1669390400
transform 1 0 21504 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0548_
timestamp 1669390400
transform 1 0 26656 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0549_
timestamp 1669390400
transform 1 0 22176 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0550_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22848 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0551_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 24192 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0552_
timestamp 1669390400
transform -1 0 26208 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0553_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 48944 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0554_
timestamp 1669390400
transform 1 0 45024 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0555_
timestamp 1669390400
transform 1 0 48944 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0556_
timestamp 1669390400
transform 1 0 49392 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0557_
timestamp 1669390400
transform 1 0 41216 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0558_
timestamp 1669390400
transform 1 0 38864 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0559_
timestamp 1669390400
transform 1 0 41440 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0560_
timestamp 1669390400
transform 1 0 41440 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0561_
timestamp 1669390400
transform 1 0 49728 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0562_
timestamp 1669390400
transform 1 0 53536 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0563_
timestamp 1669390400
transform 1 0 6720 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0564_
timestamp 1669390400
transform 1 0 5936 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0565_
timestamp 1669390400
transform -1 0 8960 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0566_
timestamp 1669390400
transform 1 0 13552 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0567_
timestamp 1669390400
transform 1 0 11760 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0568_
timestamp 1669390400
transform -1 0 18704 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0569_
timestamp 1669390400
transform -1 0 13664 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0570_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7728 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0571_
timestamp 1669390400
transform -1 0 6272 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0572_
timestamp 1669390400
transform 1 0 2576 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0573_
timestamp 1669390400
transform 1 0 12208 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0574_
timestamp 1669390400
transform -1 0 13104 0 1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0575_
timestamp 1669390400
transform 1 0 8288 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0576_
timestamp 1669390400
transform 1 0 9632 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0577_
timestamp 1669390400
transform -1 0 10640 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0578_
timestamp 1669390400
transform 1 0 12320 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0579_
timestamp 1669390400
transform 1 0 13216 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0580_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13552 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0581_
timestamp 1669390400
transform -1 0 14224 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0582_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 13216 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0583_
timestamp 1669390400
transform -1 0 11088 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0584_
timestamp 1669390400
transform -1 0 8064 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0585_
timestamp 1669390400
transform -1 0 8960 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0586_
timestamp 1669390400
transform 1 0 8288 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0587_
timestamp 1669390400
transform 1 0 7168 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0588_
timestamp 1669390400
transform -1 0 8960 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0589_
timestamp 1669390400
transform -1 0 8064 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0590_
timestamp 1669390400
transform 1 0 8288 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0591_
timestamp 1669390400
transform 1 0 9632 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0592_
timestamp 1669390400
transform -1 0 28112 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0593_
timestamp 1669390400
transform 1 0 22288 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0594_
timestamp 1669390400
transform 1 0 23296 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0595_
timestamp 1669390400
transform 1 0 24304 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0596_
timestamp 1669390400
transform -1 0 28224 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0597_
timestamp 1669390400
transform 1 0 26096 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0598_
timestamp 1669390400
transform 1 0 27104 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0599_
timestamp 1669390400
transform -1 0 28336 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0600_
timestamp 1669390400
transform -1 0 27216 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0601_
timestamp 1669390400
transform -1 0 27888 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0602_
timestamp 1669390400
transform -1 0 25088 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0603_
timestamp 1669390400
transform 1 0 21840 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0604_
timestamp 1669390400
transform -1 0 22512 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0605_
timestamp 1669390400
transform -1 0 22512 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0606_
timestamp 1669390400
transform 1 0 22736 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0607_
timestamp 1669390400
transform -1 0 23184 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0608_
timestamp 1669390400
transform -1 0 53088 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0609_
timestamp 1669390400
transform 1 0 49392 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0610_
timestamp 1669390400
transform 1 0 49392 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0611_
timestamp 1669390400
transform 1 0 51072 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0612_
timestamp 1669390400
transform 1 0 51968 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0613_
timestamp 1669390400
transform 1 0 53872 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0614_
timestamp 1669390400
transform -1 0 53648 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0615_
timestamp 1669390400
transform 1 0 53312 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0616_
timestamp 1669390400
transform -1 0 51744 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0617_
timestamp 1669390400
transform -1 0 48944 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0618_
timestamp 1669390400
transform -1 0 48832 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0619_
timestamp 1669390400
transform -1 0 48048 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0620_
timestamp 1669390400
transform 1 0 49392 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0621_
timestamp 1669390400
transform -1 0 7728 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0622_
timestamp 1669390400
transform 1 0 5824 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0623_
timestamp 1669390400
transform 1 0 5040 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0624_
timestamp 1669390400
transform 1 0 5712 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0625_
timestamp 1669390400
transform 1 0 6160 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0626_
timestamp 1669390400
transform 1 0 5936 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0627_
timestamp 1669390400
transform -1 0 6944 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0628_
timestamp 1669390400
transform 1 0 7168 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0629_
timestamp 1669390400
transform 1 0 9632 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0630_
timestamp 1669390400
transform -1 0 9184 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0631_
timestamp 1669390400
transform 1 0 38192 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0632_
timestamp 1669390400
transform -1 0 39872 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0633_
timestamp 1669390400
transform -1 0 38976 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0634_
timestamp 1669390400
transform 1 0 39200 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0635_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 40320 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0636_
timestamp 1669390400
transform -1 0 38752 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0637_
timestamp 1669390400
transform -1 0 46032 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0638_
timestamp 1669390400
transform 1 0 43456 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0639_
timestamp 1669390400
transform 1 0 45360 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0640_
timestamp 1669390400
transform 1 0 51856 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0641_
timestamp 1669390400
transform -1 0 10304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0642_
timestamp 1669390400
transform 1 0 7056 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0643_
timestamp 1669390400
transform -1 0 12656 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0644_
timestamp 1669390400
transform 1 0 14224 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _0645_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 11648 0 -1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0646_
timestamp 1669390400
transform 1 0 9744 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0647_
timestamp 1669390400
transform -1 0 6496 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0648_
timestamp 1669390400
transform 1 0 2464 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0649_
timestamp 1669390400
transform -1 0 4480 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0650_
timestamp 1669390400
transform 1 0 2800 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0651_
timestamp 1669390400
transform 1 0 9744 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0652_
timestamp 1669390400
transform 1 0 7840 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0653_
timestamp 1669390400
transform 1 0 6496 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0654_
timestamp 1669390400
transform 1 0 6496 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0655_
timestamp 1669390400
transform 1 0 8512 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0656_
timestamp 1669390400
transform -1 0 11200 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0657_
timestamp 1669390400
transform 1 0 9632 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0658_
timestamp 1669390400
transform 1 0 9632 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0659_
timestamp 1669390400
transform -1 0 11312 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0660_
timestamp 1669390400
transform 1 0 9632 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0661_
timestamp 1669390400
transform 1 0 11424 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0662_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10976 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0663_
timestamp 1669390400
transform 1 0 11984 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0664_
timestamp 1669390400
transform -1 0 13104 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0665_
timestamp 1669390400
transform 1 0 10640 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0666_
timestamp 1669390400
transform -1 0 13104 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0667_
timestamp 1669390400
transform -1 0 13104 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0668_
timestamp 1669390400
transform 1 0 10640 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0669_
timestamp 1669390400
transform -1 0 9632 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0670_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 10528 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0671_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6496 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0672_
timestamp 1669390400
transform -1 0 47376 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0673_
timestamp 1669390400
transform 1 0 46032 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0674_
timestamp 1669390400
transform -1 0 51968 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0675_
timestamp 1669390400
transform -1 0 52640 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0676_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 49392 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0677_
timestamp 1669390400
transform -1 0 48944 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0678_
timestamp 1669390400
transform 1 0 45360 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0679_
timestamp 1669390400
transform -1 0 46816 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0680_
timestamp 1669390400
transform -1 0 44912 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0681_
timestamp 1669390400
transform 1 0 45360 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0682_
timestamp 1669390400
transform -1 0 50064 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0683_
timestamp 1669390400
transform -1 0 46368 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0684_
timestamp 1669390400
transform -1 0 48384 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0685_
timestamp 1669390400
transform -1 0 48608 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0686_
timestamp 1669390400
transform -1 0 46480 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0687_
timestamp 1669390400
transform 1 0 46704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0688_
timestamp 1669390400
transform -1 0 50848 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0689_
timestamp 1669390400
transform -1 0 48944 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0690_
timestamp 1669390400
transform 1 0 52192 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0691_
timestamp 1669390400
transform 1 0 51072 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0692_
timestamp 1669390400
transform -1 0 51632 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0693_
timestamp 1669390400
transform 1 0 50736 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0694_
timestamp 1669390400
transform 1 0 52192 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0695_
timestamp 1669390400
transform -1 0 52640 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0696_
timestamp 1669390400
transform -1 0 51744 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0697_
timestamp 1669390400
transform 1 0 49392 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0698_
timestamp 1669390400
transform 1 0 51072 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0699_
timestamp 1669390400
transform -1 0 48832 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0700_
timestamp 1669390400
transform -1 0 33040 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0701_
timestamp 1669390400
transform -1 0 25088 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0702_
timestamp 1669390400
transform -1 0 31472 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0703_
timestamp 1669390400
transform -1 0 27216 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _0704_
timestamp 1669390400
transform -1 0 24640 0 1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0705_
timestamp 1669390400
transform 1 0 27328 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0706_
timestamp 1669390400
transform 1 0 28336 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0707_
timestamp 1669390400
transform -1 0 31360 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0708_
timestamp 1669390400
transform -1 0 28896 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0709_
timestamp 1669390400
transform -1 0 31248 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0710_
timestamp 1669390400
transform -1 0 32368 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0711_
timestamp 1669390400
transform 1 0 29568 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0712_
timestamp 1669390400
transform 1 0 27888 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0713_
timestamp 1669390400
transform 1 0 30576 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0714_
timestamp 1669390400
transform -1 0 30352 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0715_
timestamp 1669390400
transform -1 0 26992 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0716_
timestamp 1669390400
transform -1 0 26208 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0717_
timestamp 1669390400
transform -1 0 26432 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0718_
timestamp 1669390400
transform -1 0 26432 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0719_
timestamp 1669390400
transform -1 0 27552 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0720_
timestamp 1669390400
transform 1 0 25536 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0721_
timestamp 1669390400
transform -1 0 25088 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0722_
timestamp 1669390400
transform -1 0 26432 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0723_
timestamp 1669390400
transform 1 0 26320 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0724_
timestamp 1669390400
transform 1 0 11424 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0725_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 16800 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0726_
timestamp 1669390400
transform -1 0 16352 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0727_
timestamp 1669390400
transform 1 0 9632 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0728_
timestamp 1669390400
transform 1 0 4816 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0729_
timestamp 1669390400
transform 1 0 4032 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0730_
timestamp 1669390400
transform 1 0 6384 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0731__235 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 3808 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0731_
timestamp 1669390400
transform 1 0 1904 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0732__234
timestamp 1669390400
transform 1 0 2576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0732_
timestamp 1669390400
transform 1 0 1904 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0733__233
timestamp 1669390400
transform 1 0 16240 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0733_
timestamp 1669390400
transform -1 0 18480 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0734_
timestamp 1669390400
transform 1 0 13552 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0734__232
timestamp 1669390400
transform 1 0 13552 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0735_
timestamp 1669390400
transform 1 0 9856 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0735__231
timestamp 1669390400
transform -1 0 12096 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0736__230
timestamp 1669390400
transform -1 0 14000 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0736_
timestamp 1669390400
transform 1 0 12096 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0737__229
timestamp 1669390400
transform -1 0 16240 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0737_
timestamp 1669390400
transform 1 0 14336 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0738__228
timestamp 1669390400
transform 1 0 13664 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0738_
timestamp 1669390400
transform 1 0 13104 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0739__227
timestamp 1669390400
transform -1 0 14112 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0739_
timestamp 1669390400
transform 1 0 12656 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0740__226
timestamp 1669390400
transform 1 0 11984 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0740_
timestamp 1669390400
transform 1 0 11648 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0741__225
timestamp 1669390400
transform -1 0 6048 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0741_
timestamp 1669390400
transform 1 0 4256 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0742_
timestamp 1669390400
transform 1 0 5264 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0742__224
timestamp 1669390400
transform -1 0 6720 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0743__223
timestamp 1669390400
transform 1 0 9856 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0743_
timestamp 1669390400
transform -1 0 12208 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0744_
timestamp 1669390400
transform 1 0 5936 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0744__222
timestamp 1669390400
transform -1 0 7392 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0745_
timestamp 1669390400
transform 1 0 8176 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0745__221
timestamp 1669390400
transform -1 0 10080 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0746_
timestamp 1669390400
transform 1 0 7392 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0746__220
timestamp 1669390400
transform -1 0 8848 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0747__219
timestamp 1669390400
transform -1 0 6160 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0747_
timestamp 1669390400
transform 1 0 4704 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0748_
timestamp 1669390400
transform 1 0 5824 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0748__218
timestamp 1669390400
transform -1 0 7168 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0749__217
timestamp 1669390400
transform -1 0 7616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0749_
timestamp 1669390400
transform 1 0 6272 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0750__216
timestamp 1669390400
transform -1 0 3024 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0750_
timestamp 1669390400
transform 1 0 1680 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0751__215
timestamp 1669390400
transform -1 0 3024 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0751_
timestamp 1669390400
transform 1 0 1680 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0752_
timestamp 1669390400
transform 1 0 53424 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0753_
timestamp 1669390400
transform 1 0 22960 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0754_
timestamp 1669390400
transform -1 0 30240 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0755_
timestamp 1669390400
transform 1 0 25312 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0756_
timestamp 1669390400
transform 1 0 23856 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0757_
timestamp 1669390400
transform 1 0 18816 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0758_
timestamp 1669390400
transform 1 0 19040 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0759__214
timestamp 1669390400
transform 1 0 21616 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0759_
timestamp 1669390400
transform 1 0 21056 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0760_
timestamp 1669390400
transform 1 0 21504 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0760__213
timestamp 1669390400
transform 1 0 22064 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0761_
timestamp 1669390400
transform 1 0 17808 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0761__212
timestamp 1669390400
transform -1 0 19824 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0762__211
timestamp 1669390400
transform -1 0 25984 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0762_
timestamp 1669390400
transform 1 0 22288 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0763_
timestamp 1669390400
transform 1 0 17696 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0763__210
timestamp 1669390400
transform -1 0 19152 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0764_
timestamp 1669390400
transform 1 0 16352 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0764__209
timestamp 1669390400
transform -1 0 18032 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0765__208
timestamp 1669390400
transform -1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0765_
timestamp 1669390400
transform 1 0 19152 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0766__207
timestamp 1669390400
transform 1 0 23408 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0766_
timestamp 1669390400
transform -1 0 25760 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0767_
timestamp 1669390400
transform 1 0 25088 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0767__206
timestamp 1669390400
transform -1 0 26320 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0768__205
timestamp 1669390400
transform -1 0 24080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0768_
timestamp 1669390400
transform 1 0 21616 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0769_
timestamp 1669390400
transform 1 0 25536 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0769__204
timestamp 1669390400
transform -1 0 26768 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0770__203
timestamp 1669390400
transform -1 0 27440 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0770_
timestamp 1669390400
transform 1 0 25984 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0771__202
timestamp 1669390400
transform -1 0 30352 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0771_
timestamp 1669390400
transform 1 0 29008 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0772_
timestamp 1669390400
transform 1 0 29568 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0772__201
timestamp 1669390400
transform -1 0 31024 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0773__200
timestamp 1669390400
transform -1 0 31248 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0773_
timestamp 1669390400
transform 1 0 29792 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0774_
timestamp 1669390400
transform -1 0 36512 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0774__199
timestamp 1669390400
transform 1 0 33712 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0775_
timestamp 1669390400
transform 1 0 16688 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0775__198
timestamp 1669390400
transform -1 0 18144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0776_
timestamp 1669390400
transform 1 0 13888 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0776__197
timestamp 1669390400
transform -1 0 15904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0777__196
timestamp 1669390400
transform -1 0 17024 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0777_
timestamp 1669390400
transform 1 0 15568 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0778__195
timestamp 1669390400
transform -1 0 17024 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0778_
timestamp 1669390400
transform 1 0 15680 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0779_
timestamp 1669390400
transform 1 0 19824 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0779__194
timestamp 1669390400
transform -1 0 21952 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0780__193
timestamp 1669390400
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0780_
timestamp 1669390400
transform 1 0 20384 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0781_
timestamp 1669390400
transform -1 0 4928 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0782_
timestamp 1669390400
transform 1 0 50624 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0783_
timestamp 1669390400
transform 1 0 53312 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0784_
timestamp 1669390400
transform 1 0 49616 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0785_
timestamp 1669390400
transform 1 0 45920 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0786_
timestamp 1669390400
transform -1 0 50288 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0787__192
timestamp 1669390400
transform -1 0 35840 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0787_
timestamp 1669390400
transform 1 0 33712 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0788__191
timestamp 1669390400
transform 1 0 37408 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0788_
timestamp 1669390400
transform -1 0 40656 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0789_
timestamp 1669390400
transform 1 0 32816 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0789__190
timestamp 1669390400
transform -1 0 34160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0790__189
timestamp 1669390400
transform -1 0 33936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0790_
timestamp 1669390400
transform 1 0 31696 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0791_
timestamp 1669390400
transform 1 0 33488 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0791__188
timestamp 1669390400
transform 1 0 33824 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0792__187
timestamp 1669390400
transform 1 0 36288 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0792_
timestamp 1669390400
transform -1 0 38416 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0793_
timestamp 1669390400
transform 1 0 29008 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0793__186
timestamp 1669390400
transform -1 0 30464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0794__185
timestamp 1669390400
transform -1 0 32928 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0794_
timestamp 1669390400
transform 1 0 31360 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0795__184
timestamp 1669390400
transform 1 0 33712 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0795_
timestamp 1669390400
transform 1 0 33488 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0796__183
timestamp 1669390400
transform 1 0 34048 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0796_
timestamp 1669390400
transform 1 0 33488 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0797_
timestamp 1669390400
transform 1 0 28112 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0797__182
timestamp 1669390400
transform -1 0 29904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0798_
timestamp 1669390400
transform 1 0 29456 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0798__181
timestamp 1669390400
transform -1 0 30688 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0799__180
timestamp 1669390400
transform -1 0 29904 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0799_
timestamp 1669390400
transform 1 0 28448 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0800__179
timestamp 1669390400
transform -1 0 30464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0800_
timestamp 1669390400
transform 1 0 29120 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0801_
timestamp 1669390400
transform 1 0 40880 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0801__178
timestamp 1669390400
transform 1 0 40320 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0802_
timestamp 1669390400
transform 1 0 40768 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0802__177
timestamp 1669390400
transform -1 0 42224 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0803__176
timestamp 1669390400
transform 1 0 44352 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0803_
timestamp 1669390400
transform -1 0 45920 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0804_
timestamp 1669390400
transform -1 0 46816 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0804__175
timestamp 1669390400
transform 1 0 45360 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0805_
timestamp 1669390400
transform 1 0 39200 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0805__174
timestamp 1669390400
transform -1 0 40656 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0806_
timestamp 1669390400
transform 1 0 37744 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0806__173
timestamp 1669390400
transform -1 0 39200 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0807_
timestamp 1669390400
transform 1 0 40320 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0807__172
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0808__171
timestamp 1669390400
transform -1 0 44576 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0808_
timestamp 1669390400
transform -1 0 44912 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0809_
timestamp 1669390400
transform 1 0 31920 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0809__170
timestamp 1669390400
transform -1 0 33936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0810_
timestamp 1669390400
transform 1 0 40320 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0811_
timestamp 1669390400
transform -1 0 9184 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0812_
timestamp 1669390400
transform -1 0 6160 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0813_
timestamp 1669390400
transform 1 0 3248 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0814_
timestamp 1669390400
transform -1 0 10976 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0815__169
timestamp 1669390400
transform -1 0 23296 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0815_
timestamp 1669390400
transform 1 0 21840 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0816__168
timestamp 1669390400
transform -1 0 24976 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0816_
timestamp 1669390400
transform 1 0 23520 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0817_
timestamp 1669390400
transform 1 0 23856 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0817__167
timestamp 1669390400
transform -1 0 25088 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0818__166
timestamp 1669390400
transform 1 0 26992 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0818_
timestamp 1669390400
transform -1 0 29344 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0819__165
timestamp 1669390400
transform -1 0 23520 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0819_
timestamp 1669390400
transform 1 0 22064 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0820__164
timestamp 1669390400
transform -1 0 23632 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0820_
timestamp 1669390400
transform 1 0 21840 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0821__163
timestamp 1669390400
transform -1 0 22848 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0821_
timestamp 1669390400
transform 1 0 21392 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0822__162
timestamp 1669390400
transform 1 0 24864 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0822_
timestamp 1669390400
transform 1 0 24640 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0823_
timestamp 1669390400
transform 1 0 16128 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0823__161
timestamp 1669390400
transform -1 0 18032 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0824_
timestamp 1669390400
transform 1 0 17584 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0824__160
timestamp 1669390400
transform 1 0 18032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0825__159
timestamp 1669390400
transform -1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0825_
timestamp 1669390400
transform 1 0 18368 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0826__158
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0826_
timestamp 1669390400
transform 1 0 16464 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0827__157
timestamp 1669390400
transform -1 0 19264 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0827_
timestamp 1669390400
transform 1 0 17808 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0828__156
timestamp 1669390400
transform -1 0 18032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0828_
timestamp 1669390400
transform 1 0 15568 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0829_
timestamp 1669390400
transform 1 0 18704 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0829__155
timestamp 1669390400
transform 1 0 19264 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0830__154
timestamp 1669390400
transform 1 0 18032 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0830_
timestamp 1669390400
transform 1 0 17584 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0831__153
timestamp 1669390400
transform -1 0 11872 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0831_
timestamp 1669390400
transform 1 0 9856 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0832_
timestamp 1669390400
transform 1 0 9856 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0832__152
timestamp 1669390400
transform -1 0 11760 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0833__151
timestamp 1669390400
transform -1 0 14000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0833_
timestamp 1669390400
transform 1 0 12432 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0834__150
timestamp 1669390400
transform -1 0 14112 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0834_
timestamp 1669390400
transform 1 0 12768 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0835_
timestamp 1669390400
transform 1 0 13552 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0835__149
timestamp 1669390400
transform 1 0 13664 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0836__148
timestamp 1669390400
transform -1 0 11536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0836_
timestamp 1669390400
transform 1 0 9856 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0837__147
timestamp 1669390400
transform -1 0 14000 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0837_
timestamp 1669390400
transform 1 0 12656 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0838__146
timestamp 1669390400
transform -1 0 18032 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0838_
timestamp 1669390400
transform -1 0 17472 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0839_
timestamp 1669390400
transform 1 0 45696 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0840_
timestamp 1669390400
transform 1 0 36736 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0841_
timestamp 1669390400
transform 1 0 37408 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0842_
timestamp 1669390400
transform 1 0 37408 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0843__145
timestamp 1669390400
transform -1 0 36736 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0843_
timestamp 1669390400
transform 1 0 35392 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0844_
timestamp 1669390400
transform -1 0 41888 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0844__144
timestamp 1669390400
transform 1 0 39536 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0845_
timestamp 1669390400
transform 1 0 33488 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0845__143
timestamp 1669390400
transform 1 0 34048 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0846_
timestamp 1669390400
transform 1 0 33936 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0846__142
timestamp 1669390400
transform -1 0 35392 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0847_
timestamp 1669390400
transform 1 0 37856 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0847__141
timestamp 1669390400
transform -1 0 39200 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0848__140
timestamp 1669390400
transform -1 0 37856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0848_
timestamp 1669390400
transform 1 0 34720 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0849__139
timestamp 1669390400
transform -1 0 31920 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0849_
timestamp 1669390400
transform 1 0 29904 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0850__138
timestamp 1669390400
transform -1 0 29904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0850_
timestamp 1669390400
transform 1 0 28000 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0851_
timestamp 1669390400
transform 1 0 30464 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0851__137
timestamp 1669390400
transform -1 0 31920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0852__136
timestamp 1669390400
transform -1 0 33824 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0852_
timestamp 1669390400
transform 1 0 31808 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0853__135
timestamp 1669390400
transform -1 0 33152 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0853_
timestamp 1669390400
transform 1 0 30912 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0854_
timestamp 1669390400
transform -1 0 36736 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0854__134
timestamp 1669390400
transform 1 0 34384 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0855__133
timestamp 1669390400
transform -1 0 32704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0855_
timestamp 1669390400
transform 1 0 31248 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0856_
timestamp 1669390400
transform -1 0 35392 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0856__132
timestamp 1669390400
transform 1 0 33488 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0857__131
timestamp 1669390400
transform -1 0 28448 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0857_
timestamp 1669390400
transform 1 0 26320 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0858_
timestamp 1669390400
transform 1 0 29456 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0858__130
timestamp 1669390400
transform 1 0 29792 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0859__129
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0859_
timestamp 1669390400
transform 1 0 28336 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0860__128
timestamp 1669390400
transform -1 0 32032 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0860_
timestamp 1669390400
transform 1 0 29792 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0861__127
timestamp 1669390400
transform -1 0 25984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0861_
timestamp 1669390400
transform 1 0 23744 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0862__126
timestamp 1669390400
transform -1 0 27664 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0862_
timestamp 1669390400
transform 1 0 25760 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0863_
timestamp 1669390400
transform 1 0 27216 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0863__125
timestamp 1669390400
transform -1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0864__124
timestamp 1669390400
transform -1 0 28784 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0864_
timestamp 1669390400
transform 1 0 27440 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0865_
timestamp 1669390400
transform 1 0 29456 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0865__123
timestamp 1669390400
transform 1 0 29568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0866_
timestamp 1669390400
transform 1 0 25760 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0866__122
timestamp 1669390400
transform -1 0 27776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0867__121
timestamp 1669390400
transform -1 0 36624 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0867_
timestamp 1669390400
transform 1 0 35280 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0868_
timestamp 1669390400
transform 1 0 53200 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0869_
timestamp 1669390400
transform -1 0 46144 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0870_
timestamp 1669390400
transform -1 0 47152 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0871__120
timestamp 1669390400
transform -1 0 48384 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0871_
timestamp 1669390400
transform 1 0 47040 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0872__119
timestamp 1669390400
transform 1 0 48720 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0872_
timestamp 1669390400
transform 1 0 49392 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0873__118
timestamp 1669390400
transform 1 0 50064 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0873_
timestamp 1669390400
transform 1 0 49392 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0874_
timestamp 1669390400
transform 1 0 50960 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0874__117
timestamp 1669390400
transform -1 0 52416 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0875__116
timestamp 1669390400
transform 1 0 50400 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0875_
timestamp 1669390400
transform 1 0 49840 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0876__115
timestamp 1669390400
transform 1 0 49504 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0876_
timestamp 1669390400
transform 1 0 49392 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0877_
timestamp 1669390400
transform 1 0 51072 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0877__114
timestamp 1669390400
transform -1 0 52416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0878__113
timestamp 1669390400
transform -1 0 54320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0878_
timestamp 1669390400
transform 1 0 52864 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0879_
timestamp 1669390400
transform 1 0 43568 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0879__112
timestamp 1669390400
transform -1 0 44912 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0880__111
timestamp 1669390400
transform 1 0 45584 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0880_
timestamp 1669390400
transform 1 0 45360 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0881__110
timestamp 1669390400
transform 1 0 48160 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0881_
timestamp 1669390400
transform -1 0 52080 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0882_
timestamp 1669390400
transform 1 0 45360 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0882__109
timestamp 1669390400
transform -1 0 46704 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0883__108
timestamp 1669390400
transform 1 0 37856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0883_
timestamp 1669390400
transform 1 0 37632 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0884__107
timestamp 1669390400
transform -1 0 39984 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0884_
timestamp 1669390400
transform 1 0 38528 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0885_
timestamp 1669390400
transform 1 0 36288 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0885__106
timestamp 1669390400
transform -1 0 37856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0886__105
timestamp 1669390400
transform -1 0 42672 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0886_
timestamp 1669390400
transform 1 0 41440 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0887__104
timestamp 1669390400
transform -1 0 38640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0887_
timestamp 1669390400
transform 1 0 37408 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0888_
timestamp 1669390400
transform 1 0 35056 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0888__103
timestamp 1669390400
transform -1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0889_
timestamp 1669390400
transform 1 0 40880 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0889__102
timestamp 1669390400
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0890_
timestamp 1669390400
transform 1 0 37744 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0890__101
timestamp 1669390400
transform -1 0 39424 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0891__100
timestamp 1669390400
transform -1 0 35168 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0891_
timestamp 1669390400
transform 1 0 33824 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0892__99
timestamp 1669390400
transform 1 0 33600 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0892_
timestamp 1669390400
transform 1 0 33488 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0893__98
timestamp 1669390400
transform -1 0 35504 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0893_
timestamp 1669390400
transform 1 0 33712 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0894__97
timestamp 1669390400
transform 1 0 37408 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0894_
timestamp 1669390400
transform -1 0 40656 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0895__96
timestamp 1669390400
transform 1 0 41440 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0895_
timestamp 1669390400
transform 1 0 40880 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0896_
timestamp 1669390400
transform 1 0 39872 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0896__95
timestamp 1669390400
transform -1 0 41888 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0897_
timestamp 1669390400
transform -1 0 4928 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0898_
timestamp 1669390400
transform -1 0 53872 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0899__94
timestamp 1669390400
transform -1 0 49840 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0899_
timestamp 1669390400
transform 1 0 47936 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0900__93
timestamp 1669390400
transform -1 0 40320 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0900_
timestamp 1669390400
transform 1 0 38864 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0901_
timestamp 1669390400
transform 1 0 45360 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0901__92
timestamp 1669390400
transform 1 0 43792 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0902__91
timestamp 1669390400
transform 1 0 46032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0902_
timestamp 1669390400
transform -1 0 48608 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0903__90
timestamp 1669390400
transform 1 0 41552 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0903_
timestamp 1669390400
transform 1 0 40880 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0904__89
timestamp 1669390400
transform -1 0 43120 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0904_
timestamp 1669390400
transform 1 0 41664 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0905_
timestamp 1669390400
transform 1 0 42336 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0905__88
timestamp 1669390400
transform -1 0 45808 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0906__87
timestamp 1669390400
transform 1 0 46368 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0906_
timestamp 1669390400
transform -1 0 48608 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0907_
timestamp 1669390400
transform -1 0 48608 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0907__86
timestamp 1669390400
transform 1 0 43792 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0908_
timestamp 1669390400
transform 1 0 41440 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0908__85
timestamp 1669390400
transform 1 0 40768 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0909__84
timestamp 1669390400
transform -1 0 44016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0909_
timestamp 1669390400
transform 1 0 42560 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0910__83
timestamp 1669390400
transform 1 0 46256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0910_
timestamp 1669390400
transform -1 0 48608 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0911__82
timestamp 1669390400
transform 1 0 48944 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0911_
timestamp 1669390400
transform 1 0 49392 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0912__81
timestamp 1669390400
transform -1 0 48720 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0912_
timestamp 1669390400
transform 1 0 47264 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0913__80
timestamp 1669390400
transform -1 0 53760 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0913_
timestamp 1669390400
transform 1 0 49616 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0914__79
timestamp 1669390400
transform 1 0 53872 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0914_
timestamp 1669390400
transform -1 0 56560 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0915__78
timestamp 1669390400
transform -1 0 50848 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0915_
timestamp 1669390400
transform 1 0 48720 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0916__77
timestamp 1669390400
transform 1 0 49728 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0916_
timestamp 1669390400
transform 1 0 49392 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0917_
timestamp 1669390400
transform -1 0 56560 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0917__76
timestamp 1669390400
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0918__75
timestamp 1669390400
transform 1 0 54544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0918_
timestamp 1669390400
transform -1 0 56896 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0919__74
timestamp 1669390400
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0919_
timestamp 1669390400
transform 1 0 48832 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0920__73
timestamp 1669390400
transform -1 0 47488 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0920_
timestamp 1669390400
transform 1 0 46032 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0921__72
timestamp 1669390400
transform 1 0 50176 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0921_
timestamp 1669390400
transform 1 0 49504 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0922__71
timestamp 1669390400
transform -1 0 55664 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0922_
timestamp 1669390400
transform -1 0 55440 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0923__70
timestamp 1669390400
transform 1 0 48384 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0923_
timestamp 1669390400
transform 1 0 49392 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0924__69
timestamp 1669390400
transform 1 0 54656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0924_
timestamp 1669390400
transform -1 0 56560 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0925__68
timestamp 1669390400
transform 1 0 42000 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0925_
timestamp 1669390400
transform 1 0 41440 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0926_
timestamp 1669390400
transform 1 0 53648 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0927_
timestamp 1669390400
transform 1 0 1904 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0928_
timestamp 1669390400
transform 1 0 1680 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0929_
timestamp 1669390400
transform 1 0 5600 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0930_
timestamp 1669390400
transform 1 0 5600 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0931_
timestamp 1669390400
transform 1 0 8288 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0932_
timestamp 1669390400
transform -1 0 15680 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0933_
timestamp 1669390400
transform 1 0 12544 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0934_
timestamp 1669390400
transform 1 0 10752 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0935_
timestamp 1669390400
transform 1 0 7728 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0936_
timestamp 1669390400
transform 1 0 3248 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0937__67
timestamp 1669390400
transform -1 0 10080 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0937_
timestamp 1669390400
transform 1 0 8512 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0938_
timestamp 1669390400
transform 1 0 9520 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0938__66
timestamp 1669390400
transform -1 0 10976 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0939_
timestamp 1669390400
transform 1 0 11200 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0939__65
timestamp 1669390400
transform -1 0 12544 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0940__64
timestamp 1669390400
transform 1 0 14672 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0940_
timestamp 1669390400
transform -1 0 16240 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0941_
timestamp 1669390400
transform 1 0 5936 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0941__63
timestamp 1669390400
transform -1 0 7616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0942_
timestamp 1669390400
transform 1 0 9632 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0942__62
timestamp 1669390400
transform -1 0 10976 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0943_
timestamp 1669390400
transform 1 0 8848 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0943__61
timestamp 1669390400
transform -1 0 10192 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0944_
timestamp 1669390400
transform 1 0 9184 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0944__60
timestamp 1669390400
transform -1 0 10640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0945__59
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0945_
timestamp 1669390400
transform 1 0 13552 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0946__58
timestamp 1669390400
transform -1 0 15120 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0946_
timestamp 1669390400
transform 1 0 13776 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0947__57
timestamp 1669390400
transform -1 0 16352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0947_
timestamp 1669390400
transform 1 0 14336 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0948__56
timestamp 1669390400
transform -1 0 15792 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0948_
timestamp 1669390400
transform 1 0 13888 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0949__55
timestamp 1669390400
transform -1 0 6832 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0949_
timestamp 1669390400
transform 1 0 5488 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0950__54
timestamp 1669390400
transform -1 0 4928 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0950_
timestamp 1669390400
transform 1 0 2464 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0951__53
timestamp 1669390400
transform -1 0 3472 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0951_
timestamp 1669390400
transform 1 0 2016 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0952__52
timestamp 1669390400
transform -1 0 4144 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0952_
timestamp 1669390400
transform 1 0 1904 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0953_
timestamp 1669390400
transform -1 0 5264 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0953__51
timestamp 1669390400
transform -1 0 4816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0954__50
timestamp 1669390400
transform -1 0 6832 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0954_
timestamp 1669390400
transform 1 0 5488 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0955_
timestamp 1669390400
transform 1 0 24192 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0956_
timestamp 1669390400
transform 1 0 41664 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0957_
timestamp 1669390400
transform 1 0 43344 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0958_
timestamp 1669390400
transform 1 0 42000 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0959_
timestamp 1669390400
transform -1 0 48272 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0960_
timestamp 1669390400
transform 1 0 47824 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0961_
timestamp 1669390400
transform -1 0 54656 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0962_
timestamp 1669390400
transform -1 0 55552 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0963_
timestamp 1669390400
transform 1 0 49616 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0964_
timestamp 1669390400
transform 1 0 46256 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0965__49
timestamp 1669390400
transform -1 0 39984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0965_
timestamp 1669390400
transform 1 0 37744 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0966_
timestamp 1669390400
transform 1 0 39088 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0966__48
timestamp 1669390400
transform -1 0 40880 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0967_
timestamp 1669390400
transform 1 0 33488 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0967__47
timestamp 1669390400
transform 1 0 34160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0968__46
timestamp 1669390400
transform -1 0 36624 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0968_
timestamp 1669390400
transform 1 0 35168 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0969__45
timestamp 1669390400
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0969_
timestamp 1669390400
transform 1 0 36960 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0970__44
timestamp 1669390400
transform 1 0 37744 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0970_
timestamp 1669390400
transform 1 0 37408 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0971__43
timestamp 1669390400
transform 1 0 37408 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0971_
timestamp 1669390400
transform 1 0 37408 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0972__42
timestamp 1669390400
transform -1 0 38528 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0972_
timestamp 1669390400
transform 1 0 36064 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0973__41
timestamp 1669390400
transform -1 0 39200 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0973_
timestamp 1669390400
transform 1 0 37744 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0974__40
timestamp 1669390400
transform -1 0 41888 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0974_
timestamp 1669390400
transform 1 0 39872 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0975_
timestamp 1669390400
transform 1 0 41440 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0975__39
timestamp 1669390400
transform -1 0 43792 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0976_
timestamp 1669390400
transform 1 0 41440 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0976__38
timestamp 1669390400
transform 1 0 42000 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0977_
timestamp 1669390400
transform 1 0 42672 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0977__37
timestamp 1669390400
transform -1 0 44128 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0978__36
timestamp 1669390400
transform -1 0 44576 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0978_
timestamp 1669390400
transform 1 0 43232 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0979_
timestamp 1669390400
transform 1 0 45920 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0979__35
timestamp 1669390400
transform -1 0 48048 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0980__34
timestamp 1669390400
transform -1 0 47152 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0980_
timestamp 1669390400
transform 1 0 45696 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0981_
timestamp 1669390400
transform 1 0 45472 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0981__33
timestamp 1669390400
transform -1 0 46816 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0982__32
timestamp 1669390400
transform 1 0 49616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0982_
timestamp 1669390400
transform 1 0 49392 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0983__31
timestamp 1669390400
transform -1 0 41328 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0983_
timestamp 1669390400
transform 1 0 37744 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0984_
timestamp 1669390400
transform -1 0 5152 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0985_
timestamp 1669390400
transform 1 0 28224 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0986_
timestamp 1669390400
transform 1 0 27440 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0987_
timestamp 1669390400
transform -1 0 33936 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0988_
timestamp 1669390400
transform 1 0 27664 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0989_
timestamp 1669390400
transform -1 0 26656 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0990_
timestamp 1669390400
transform 1 0 21616 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0991_
timestamp 1669390400
transform 1 0 24864 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0992_
timestamp 1669390400
transform -1 0 26096 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0993_
timestamp 1669390400
transform 1 0 16912 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0993__30
timestamp 1669390400
transform -1 0 18256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0994_
timestamp 1669390400
transform 1 0 17584 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0994__29
timestamp 1669390400
transform 1 0 17808 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0995__28
timestamp 1669390400
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0995_
timestamp 1669390400
transform 1 0 20048 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0996__27
timestamp 1669390400
transform -1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0996_
timestamp 1669390400
transform 1 0 19264 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0997_
timestamp 1669390400
transform 1 0 24416 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0997__26
timestamp 1669390400
transform -1 0 25984 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0998__25
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0998_
timestamp 1669390400
transform 1 0 24416 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _0999__24
timestamp 1669390400
transform 1 0 26768 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _0999_
timestamp 1669390400
transform -1 0 28784 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1000__23
timestamp 1669390400
transform -1 0 24640 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1000_
timestamp 1669390400
transform 1 0 22064 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1001_
timestamp 1669390400
transform 1 0 17808 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1001__22
timestamp 1669390400
transform -1 0 20048 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1002__21
timestamp 1669390400
transform -1 0 19152 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1002_
timestamp 1669390400
transform 1 0 17696 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1003__20
timestamp 1669390400
transform -1 0 22288 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1003_
timestamp 1669390400
transform 1 0 20944 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1004_
timestamp 1669390400
transform 1 0 19488 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1004__19
timestamp 1669390400
transform -1 0 21952 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1005__18
timestamp 1669390400
transform -1 0 21952 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1005_
timestamp 1669390400
transform 1 0 19824 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1006__17
timestamp 1669390400
transform -1 0 19824 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1006_
timestamp 1669390400
transform 1 0 18368 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1007__16
timestamp 1669390400
transform -1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1007_
timestamp 1669390400
transform 1 0 14224 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1008_
timestamp 1669390400
transform 1 0 17696 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1008__15
timestamp 1669390400
transform -1 0 19040 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1009__14
timestamp 1669390400
transform -1 0 19824 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1009_
timestamp 1669390400
transform 1 0 17808 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1010_
timestamp 1669390400
transform 1 0 14336 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1010__13
timestamp 1669390400
transform -1 0 18032 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1011__12
timestamp 1669390400
transform -1 0 19600 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1011_
timestamp 1669390400
transform 1 0 18144 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  _1012__11
timestamp 1669390400
transform -1 0 21056 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1012_
timestamp 1669390400
transform 1 0 19712 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1013_
timestamp 1669390400
transform 1 0 18928 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1014_
timestamp 1669390400
transform 1 0 9856 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 29792 0 1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1669390400
transform 1 0 15232 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1669390400
transform -1 0 17024 0 -1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1669390400
transform 1 0 41776 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1669390400
transform 1 0 41776 0 -1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_0_clk
timestamp 1669390400
transform -1 0 9184 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_1_clk
timestamp 1669390400
transform 1 0 7504 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_2_clk
timestamp 1669390400
transform 1 0 5600 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_3_clk
timestamp 1669390400
transform 1 0 11424 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_4_clk
timestamp 1669390400
transform 1 0 17584 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_5_clk
timestamp 1669390400
transform 1 0 25536 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_6_clk
timestamp 1669390400
transform 1 0 18928 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_7_clk
timestamp 1669390400
transform 1 0 14112 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_8_clk
timestamp 1669390400
transform -1 0 15232 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_9_clk
timestamp 1669390400
transform 1 0 6832 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_10_clk
timestamp 1669390400
transform -1 0 15568 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_11_clk
timestamp 1669390400
transform -1 0 8848 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_12_clk
timestamp 1669390400
transform -1 0 9184 0 -1 51744
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_13_clk
timestamp 1669390400
transform 1 0 13552 0 1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_14_clk
timestamp 1669390400
transform 1 0 18256 0 -1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_15_clk
timestamp 1669390400
transform 1 0 26544 0 -1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_16_clk
timestamp 1669390400
transform 1 0 27104 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_17_clk
timestamp 1669390400
transform 1 0 19488 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_18_clk
timestamp 1669390400
transform 1 0 25536 0 -1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_19_clk
timestamp 1669390400
transform -1 0 36512 0 1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_20_clk
timestamp 1669390400
transform 1 0 34384 0 -1 39200
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_21_clk
timestamp 1669390400
transform -1 0 44128 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_22_clk
timestamp 1669390400
transform 1 0 33600 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_23_clk
timestamp 1669390400
transform 1 0 35392 0 -1 50176
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_24_clk
timestamp 1669390400
transform 1 0 42000 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_25_clk
timestamp 1669390400
transform 1 0 49392 0 -1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_26_clk
timestamp 1669390400
transform 1 0 51072 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_27_clk
timestamp 1669390400
transform -1 0 52864 0 1 39200
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_29_clk
timestamp 1669390400
transform -1 0 52864 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_30_clk
timestamp 1669390400
transform 1 0 42224 0 -1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_31_clk
timestamp 1669390400
transform 1 0 37520 0 1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_32_clk
timestamp 1669390400
transform -1 0 40992 0 -1 26656
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_33_clk
timestamp 1669390400
transform 1 0 41440 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_34_clk
timestamp 1669390400
transform 1 0 49392 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_35_clk
timestamp 1669390400
transform 1 0 51296 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_36_clk
timestamp 1669390400
transform 1 0 49392 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_37_clk
timestamp 1669390400
transform 1 0 51296 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_38_clk
timestamp 1669390400
transform 1 0 49392 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_39_clk
timestamp 1669390400
transform -1 0 47600 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_40_clk
timestamp 1669390400
transform -1 0 44912 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_41_clk
timestamp 1669390400
transform -1 0 35952 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_42_clk
timestamp 1669390400
transform 1 0 37968 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_43_clk
timestamp 1669390400
transform 1 0 33488 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_44_clk
timestamp 1669390400
transform 1 0 26768 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_45_clk
timestamp 1669390400
transform 1 0 23408 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_46_clk
timestamp 1669390400
transform 1 0 19264 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_47_clk
timestamp 1669390400
transform 1 0 26544 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_48_clk
timestamp 1669390400
transform 1 0 19488 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_49_clk
timestamp 1669390400
transform 1 0 14560 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_50_clk
timestamp 1669390400
transform -1 0 9184 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 56336 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output2
timestamp 1669390400
transform 1 0 1680 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output3
timestamp 1669390400
transform 1 0 49168 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output4
timestamp 1669390400
transform 1 0 44800 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output5
timestamp 1669390400
transform 1 0 1680 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output6
timestamp 1669390400
transform -1 0 56336 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output7
timestamp 1669390400
transform 1 0 21616 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output8
timestamp 1669390400
transform 1 0 5600 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output9
timestamp 1669390400
transform 1 0 26992 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output10
timestamp 1669390400
transform -1 0 56336 0 -1 26656
box -86 -86 1654 870
<< labels >>
flabel metal3 s 200 43680 800 43792 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 59200 5376 59800 5488 0 FreeSans 448 0 0 0 cout1
port 1 nsew signal tristate
flabel metal2 s 0 200 112 800 0 FreeSans 448 90 0 0 cout10
port 2 nsew signal tristate
flabel metal2 s 49056 59200 49168 59800 0 FreeSans 448 90 0 0 cout2
port 3 nsew signal tristate
flabel metal2 s 43680 200 43792 800 0 FreeSans 448 90 0 0 cout3
port 4 nsew signal tristate
flabel metal3 s 200 21504 800 21616 0 FreeSans 448 0 0 0 cout4
port 5 nsew signal tristate
flabel metal3 s 59200 49056 59800 49168 0 FreeSans 448 0 0 0 cout5
port 6 nsew signal tristate
flabel metal2 s 21504 200 21616 800 0 FreeSans 448 90 0 0 cout6
port 7 nsew signal tristate
flabel metal2 s 5376 59200 5488 59800 0 FreeSans 448 90 0 0 cout7
port 8 nsew signal tristate
flabel metal2 s 26880 59200 26992 59800 0 FreeSans 448 90 0 0 cout8
port 9 nsew signal tristate
flabel metal3 s 59200 26880 59800 26992 0 FreeSans 448 0 0 0 cout9
port 10 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 11 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 12 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 12 nsew ground bidirectional
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal3 3416 5992 3416 5992 0 _0000_
rlabel metal2 54152 6552 54152 6552 0 _0001_
rlabel metal3 47152 50008 47152 50008 0 _0002_
rlabel metal3 40712 5208 40712 5208 0 _0003_
rlabel metal2 3976 22960 3976 22960 0 _0004_
rlabel metal2 54376 47768 54376 47768 0 _0005_
rlabel metal2 19768 5992 19768 5992 0 _0006_
rlabel metal2 4200 51296 4200 51296 0 _0007_
rlabel metal3 25424 49672 25424 49672 0 _0008_
rlabel metal2 54040 26684 54040 26684 0 _0009_
rlabel metal2 13944 50176 13944 50176 0 _0010_
rlabel metal2 13720 45752 13720 45752 0 _0011_
rlabel metal2 10584 46312 10584 46312 0 _0012_
rlabel metal3 7392 46760 7392 46760 0 _0013_
rlabel metal3 6160 48328 6160 48328 0 _0014_
rlabel metal2 7336 50232 7336 50232 0 _0015_
rlabel metal2 23912 6832 23912 6832 0 _0037_
rlabel metal2 27832 7000 27832 7000 0 _0038_
rlabel metal2 26488 11256 26488 11256 0 _0039_
rlabel metal2 24808 8960 24808 8960 0 _0040_
rlabel metal2 21840 8456 21840 8456 0 _0041_
rlabel metal3 21336 7336 21336 7336 0 _0042_
rlabel metal2 51352 39648 51352 39648 0 _0065_
rlabel metal3 53592 38584 53592 38584 0 _0066_
rlabel metal2 50568 36792 50568 36792 0 _0067_
rlabel metal2 46928 36344 46928 36344 0 _0068_
rlabel metal2 49336 38584 49336 38584 0 _0069_
rlabel metal2 7448 29008 7448 29008 0 _0093_
rlabel metal2 5208 30632 5208 30632 0 _0094_
rlabel metal3 5208 26152 5208 26152 0 _0095_
rlabel metal2 10024 25704 10024 25704 0 _0096_
rlabel metal2 38472 11760 38472 11760 0 _0121_
rlabel metal2 38416 9912 38416 9912 0 _0122_
rlabel metal2 38360 7056 38360 7056 0 _0123_
rlabel metal2 45192 47152 45192 47152 0 _0149_
rlabel metal2 45864 49280 45864 49280 0 _0150_
rlabel metal2 52360 11816 52360 11816 0 _0177_
rlabel metal2 2856 7896 2856 7896 0 _0205_
rlabel metal2 2632 9968 2632 9968 0 _0206_
rlabel metal3 6664 11256 6664 11256 0 _0207_
rlabel metal3 8344 8344 8344 8344 0 _0208_
rlabel metal2 9240 7056 9240 7056 0 _0209_
rlabel metal3 13440 7560 13440 7560 0 _0210_
rlabel metal3 12264 9128 12264 9128 0 _0211_
rlabel metal2 11704 12488 11704 12488 0 _0212_
rlabel metal2 9240 13552 9240 13552 0 _0213_
rlabel metal3 5600 13048 5600 13048 0 _0214_
rlabel metal2 42616 24304 42616 24304 0 _0233_
rlabel metal2 44352 25704 44352 25704 0 _0234_
rlabel metal2 47656 21896 47656 21896 0 _0235_
rlabel metal2 47376 20104 47376 20104 0 _0236_
rlabel metal2 48720 20888 48720 20888 0 _0237_
rlabel metal3 52864 21224 52864 21224 0 _0238_
rlabel metal3 53648 24136 53648 24136 0 _0239_
rlabel metal2 50960 28504 50960 28504 0 _0240_
rlabel metal2 48440 26712 48440 26712 0 _0241_
rlabel metal2 29176 47152 29176 47152 0 _0261_
rlabel metal2 28392 49448 28392 49448 0 _0262_
rlabel metal3 31416 45640 31416 45640 0 _0263_
rlabel metal2 28616 43680 28616 43680 0 _0264_
rlabel metal2 25704 42224 25704 42224 0 _0265_
rlabel metal3 24696 44184 24696 44184 0 _0266_
rlabel metal2 25760 46760 25760 46760 0 _0267_
rlabel metal3 25872 48888 25872 48888 0 _0268_
rlabel metal3 11256 50008 11256 50008 0 _0289_
rlabel metal3 29736 47432 29736 47432 0 _0290_
rlabel metal3 24528 49560 24528 49560 0 _0291_
rlabel metal2 25592 45528 25592 45528 0 _0292_
rlabel metal2 25704 47824 25704 47824 0 _0293_
rlabel metal3 25424 45304 25424 45304 0 _0294_
rlabel metal3 26208 42168 26208 42168 0 _0295_
rlabel metal3 29400 48888 29400 48888 0 _0296_
rlabel metal2 30240 46088 30240 46088 0 _0297_
rlabel metal2 29848 46648 29848 46648 0 _0298_
rlabel metal2 25928 44688 25928 44688 0 _0299_
rlabel metal3 30520 44296 30520 44296 0 _0300_
rlabel metal2 26040 42672 26040 42672 0 _0301_
rlabel metal3 25200 44520 25200 44520 0 _0302_
rlabel metal2 26152 44744 26152 44744 0 _0303_
rlabel metal2 26040 47320 26040 47320 0 _0304_
rlabel metal3 25480 46536 25480 46536 0 _0305_
rlabel metal2 53368 12936 53368 12936 0 _0306_
rlabel metal2 53704 13440 53704 13440 0 _0307_
rlabel metal2 54264 8008 54264 8008 0 _0308_
rlabel metal2 54208 11592 54208 11592 0 _0309_
rlabel metal3 52808 12712 52808 12712 0 _0310_
rlabel metal3 46928 11256 46928 11256 0 _0311_
rlabel metal3 46592 11144 46592 11144 0 _0312_
rlabel metal2 46872 13216 46872 13216 0 _0313_
rlabel metal3 49784 11368 49784 11368 0 _0314_
rlabel metal2 48440 46704 48440 46704 0 _0315_
rlabel metal3 52136 46536 52136 46536 0 _0316_
rlabel metal2 48552 45584 48552 45584 0 _0317_
rlabel metal2 41608 46872 41608 46872 0 _0318_
rlabel metal2 41720 46872 41720 46872 0 _0319_
rlabel metal2 42392 45416 42392 45416 0 _0320_
rlabel metal3 42560 46648 42560 46648 0 _0321_
rlabel metal2 47096 46536 47096 46536 0 _0322_
rlabel metal2 45864 47264 45864 47264 0 _0323_
rlabel metal2 37632 16856 37632 16856 0 _0324_
rlabel metal2 38248 17696 38248 17696 0 _0325_
rlabel metal2 37352 17024 37352 17024 0 _0326_
rlabel metal2 31416 22036 31416 22036 0 _0327_
rlabel metal3 30968 23800 30968 23800 0 _0328_
rlabel metal2 31752 24808 31752 24808 0 _0329_
rlabel metal3 33264 23912 33264 23912 0 _0330_
rlabel metal3 34608 23576 34608 23576 0 _0331_
rlabel metal2 39536 5992 39536 5992 0 _0332_
rlabel metal2 15232 27608 15232 27608 0 _0333_
rlabel metal2 15568 28392 15568 28392 0 _0334_
rlabel metal2 20776 28952 20776 28952 0 _0335_
rlabel metal2 20888 26824 20888 26824 0 _0336_
rlabel metal2 21224 28168 21224 28168 0 _0337_
rlabel metal2 21560 27888 21560 27888 0 _0338_
rlabel metal2 15736 28280 15736 28280 0 _0339_
rlabel metal2 9464 27776 9464 27776 0 _0340_
rlabel metal3 7112 28840 7112 28840 0 _0341_
rlabel metal3 43736 39032 43736 39032 0 _0342_
rlabel metal2 43120 38808 43120 38808 0 _0343_
rlabel metal2 35672 40600 35672 40600 0 _0344_
rlabel metal2 37464 37240 37464 37240 0 _0345_
rlabel metal2 36568 32984 36568 32984 0 _0346_
rlabel metal3 37352 37912 37352 37912 0 _0347_
rlabel metal3 40656 37464 40656 37464 0 _0348_
rlabel metal2 48216 37968 48216 37968 0 _0349_
rlabel metal2 53032 39144 53032 39144 0 _0350_
rlabel metal3 21672 13048 21672 13048 0 _0351_
rlabel metal2 23912 12544 23912 12544 0 _0352_
rlabel metal2 28616 12488 28616 12488 0 _0353_
rlabel metal2 32200 11368 32200 11368 0 _0354_
rlabel metal3 26096 12152 26096 12152 0 _0355_
rlabel metal2 23352 17528 23352 17528 0 _0356_
rlabel metal2 23576 17864 23576 17864 0 _0357_
rlabel metal2 23688 11704 23688 11704 0 _0358_
rlabel metal3 23184 8232 23184 8232 0 _0359_
rlabel metal2 6160 41720 6160 41720 0 _0360_
rlabel metal2 9912 44632 9912 44632 0 _0361_
rlabel metal3 15232 42728 15232 42728 0 _0362_
rlabel metal3 15344 42952 15344 42952 0 _0363_
rlabel metal2 10192 44296 10192 44296 0 _0364_
rlabel metal2 8680 37408 8680 37408 0 _0365_
rlabel metal3 10192 44296 10192 44296 0 _0366_
rlabel metal2 9016 48384 9016 48384 0 _0367_
rlabel metal2 22232 48160 22232 48160 0 _0368_
rlabel metal2 22008 46984 22008 46984 0 _0369_
rlabel metal2 23240 47880 23240 47880 0 _0370_
rlabel metal2 22568 41048 22568 41048 0 _0371_
rlabel metal2 26936 40040 26936 40040 0 _0372_
rlabel metal2 23240 35112 23240 35112 0 _0373_
rlabel metal2 23464 47208 23464 47208 0 _0374_
rlabel metal3 25368 48440 25368 48440 0 _0375_
rlabel metal2 48496 26264 48496 26264 0 _0376_
rlabel metal3 47768 29288 47768 29288 0 _0377_
rlabel metal2 49728 29400 49728 29400 0 _0378_
rlabel metal2 50120 28112 50120 28112 0 _0379_
rlabel metal2 41832 22568 41832 22568 0 _0380_
rlabel metal3 40824 27048 40824 27048 0 _0381_
rlabel metal2 42056 26488 42056 26488 0 _0382_
rlabel metal3 48720 26376 48720 26376 0 _0383_
rlabel metal2 53704 26600 53704 26600 0 _0384_
rlabel metal2 7560 13832 7560 13832 0 _0385_
rlabel metal2 7224 18704 7224 18704 0 _0386_
rlabel metal2 8568 13832 8568 13832 0 _0387_
rlabel metal2 13496 17136 13496 17136 0 _0388_
rlabel metal2 12768 22232 12768 22232 0 _0389_
rlabel metal2 13160 18312 13160 18312 0 _0390_
rlabel metal3 11536 13720 11536 13720 0 _0391_
rlabel metal3 6944 12936 6944 12936 0 _0392_
rlabel metal3 3472 6664 3472 6664 0 _0393_
rlabel metal2 13160 48496 13160 48496 0 _0394_
rlabel metal2 7672 47320 7672 47320 0 _0395_
rlabel metal2 9800 46200 9800 46200 0 _0396_
rlabel metal2 10640 45864 10640 45864 0 _0397_
rlabel metal2 13608 48944 13608 48944 0 _0398_
rlabel metal2 13384 49728 13384 49728 0 _0399_
rlabel metal2 14168 45192 14168 45192 0 _0400_
rlabel metal2 10808 47096 10808 47096 0 _0401_
rlabel metal2 8344 47880 8344 47880 0 _0402_
rlabel metal2 8568 47376 8568 47376 0 _0403_
rlabel metal2 7784 48216 7784 48216 0 _0404_
rlabel metal2 7784 48048 7784 48048 0 _0405_
rlabel metal3 9296 49896 9296 49896 0 _0406_
rlabel metal2 24696 9520 24696 9520 0 _0407_
rlabel metal3 23856 10472 23856 10472 0 _0408_
rlabel metal2 22792 7168 22792 7168 0 _0409_
rlabel metal2 27496 7448 27496 7448 0 _0410_
rlabel metal3 26936 6664 26936 6664 0 _0411_
rlabel metal2 27048 11312 27048 11312 0 _0412_
rlabel metal3 26264 9800 26264 9800 0 _0413_
rlabel metal2 22904 9016 22904 9016 0 _0414_
rlabel metal2 22288 10024 22288 10024 0 _0415_
rlabel metal2 23016 7784 23016 7784 0 _0416_
rlabel metal2 49784 37912 49784 37912 0 _0417_
rlabel metal2 50120 38136 50120 38136 0 _0418_
rlabel metal2 49784 38976 49784 38976 0 _0419_
rlabel metal2 53256 37968 53256 37968 0 _0420_
rlabel metal3 53760 38696 53760 38696 0 _0421_
rlabel metal3 52584 37240 52584 37240 0 _0422_
rlabel metal2 48552 37968 48552 37968 0 _0423_
rlabel metal3 48664 38808 48664 38808 0 _0424_
rlabel metal2 6552 28896 6552 28896 0 _0425_
rlabel metal2 5544 29736 5544 29736 0 _0426_
rlabel metal2 7560 26544 7560 26544 0 _0427_
rlabel metal2 6664 26376 6664 26376 0 _0428_
rlabel metal3 8344 26040 8344 26040 0 _0429_
rlabel metal2 9464 26264 9464 26264 0 _0430_
rlabel metal2 38696 9632 38696 9632 0 _0431_
rlabel metal2 39424 10360 39424 10360 0 _0432_
rlabel metal3 38864 7336 38864 7336 0 _0433_
rlabel metal3 45136 48888 45136 48888 0 _0434_
rlabel metal2 10920 13832 10920 13832 0 _0435_
rlabel metal2 8232 9912 8232 9912 0 _0436_
rlabel metal2 11872 8232 11872 8232 0 _0437_
rlabel metal3 12208 11928 12208 11928 0 _0438_
rlabel metal2 11368 8316 11368 8316 0 _0439_
rlabel metal3 3192 7448 3192 7448 0 _0440_
rlabel metal2 3192 7980 3192 7980 0 _0441_
rlabel metal2 3416 10472 3416 10472 0 _0442_
rlabel metal2 6888 12488 6888 12488 0 _0443_
rlabel metal3 7672 9912 7672 9912 0 _0444_
rlabel metal2 7448 10080 7448 10080 0 _0445_
rlabel metal3 9632 8792 9632 8792 0 _0446_
rlabel metal3 11144 7336 11144 7336 0 _0447_
rlabel metal2 11032 8176 11032 8176 0 _0448_
rlabel metal2 10248 7728 10248 7728 0 _0449_
rlabel metal2 11760 6104 11760 6104 0 _0450_
rlabel metal2 12264 10136 12264 10136 0 _0451_
rlabel metal3 11648 9688 11648 9688 0 _0452_
rlabel metal2 12824 12264 12824 12264 0 _0453_
rlabel metal3 11648 12824 11648 12824 0 _0454_
rlabel metal2 7224 12544 7224 12544 0 _0455_
rlabel metal2 45864 23576 45864 23576 0 _0456_
rlabel metal2 48328 23240 48328 23240 0 _0457_
rlabel metal2 51128 25872 51128 25872 0 _0458_
rlabel metal3 50232 25368 50232 25368 0 _0459_
rlabel via2 49896 25480 49896 25480 0 _0460_
rlabel metal2 45472 24808 45472 24808 0 _0461_
rlabel metal3 45136 25368 45136 25368 0 _0462_
rlabel metal2 47768 23016 47768 23016 0 _0463_
rlabel metal3 47544 22344 47544 22344 0 _0464_
rlabel metal2 46088 21840 46088 21840 0 _0465_
rlabel metal2 48104 23184 48104 23184 0 _0466_
rlabel metal2 46312 20888 46312 20888 0 _0467_
rlabel metal2 49168 23128 49168 23128 0 _0468_
rlabel metal2 52024 22512 52024 22512 0 _0469_
rlabel metal2 51408 26040 51408 26040 0 _0470_
rlabel metal2 52360 24360 52360 24360 0 _0471_
rlabel metal3 51968 26936 51968 26936 0 _0472_
rlabel metal2 51352 24808 51352 24808 0 _0473_
rlabel metal2 50176 25704 50176 25704 0 _0474_
rlabel metal3 2478 43736 2478 43736 0 clk
rlabel metal2 15456 28616 15456 28616 0 clknet_0_clk
rlabel metal2 6664 22680 6664 22680 0 clknet_2_0__leaf_clk
rlabel metal2 8344 43456 8344 43456 0 clknet_2_1__leaf_clk
rlabel metal2 47320 22680 47320 22680 0 clknet_2_2__leaf_clk
rlabel metal3 46144 31752 46144 31752 0 clknet_2_3__leaf_clk
rlabel metal3 2968 12040 2968 12040 0 clknet_leaf_0_clk
rlabel metal2 6104 42336 6104 42336 0 clknet_leaf_10_clk
rlabel metal2 1960 45080 1960 45080 0 clknet_leaf_11_clk
rlabel metal2 4984 50904 4984 50904 0 clknet_leaf_12_clk
rlabel metal2 13272 50904 13272 50904 0 clknet_leaf_13_clk
rlabel metal2 22904 46256 22904 46256 0 clknet_leaf_14_clk
rlabel metal2 25928 49728 25928 49728 0 clknet_leaf_15_clk
rlabel metal2 26488 42336 26488 42336 0 clknet_leaf_16_clk
rlabel metal3 21336 44296 21336 44296 0 clknet_leaf_17_clk
rlabel metal2 24584 38808 24584 38808 0 clknet_leaf_18_clk
rlabel metal2 29960 30184 29960 30184 0 clknet_leaf_19_clk
rlabel metal2 8008 14784 8008 14784 0 clknet_leaf_1_clk
rlabel metal3 33040 37240 33040 37240 0 clknet_leaf_20_clk
rlabel metal2 40936 40320 40936 40320 0 clknet_leaf_21_clk
rlabel metal2 33656 41216 33656 41216 0 clknet_leaf_22_clk
rlabel metal3 35168 50456 35168 50456 0 clknet_leaf_23_clk
rlabel metal2 44408 45360 44408 45360 0 clknet_leaf_24_clk
rlabel metal2 45864 46256 45864 46256 0 clknet_leaf_25_clk
rlabel metal2 52696 44744 52696 44744 0 clknet_leaf_26_clk
rlabel metal3 47152 39704 47152 39704 0 clknet_leaf_27_clk
rlabel metal2 49560 31304 49560 31304 0 clknet_leaf_29_clk
rlabel metal3 3976 21896 3976 21896 0 clknet_leaf_2_clk
rlabel metal3 45584 32424 45584 32424 0 clknet_leaf_30_clk
rlabel metal3 35392 29400 35392 29400 0 clknet_leaf_31_clk
rlabel metal2 35112 27440 35112 27440 0 clknet_leaf_32_clk
rlabel metal3 45920 24920 45920 24920 0 clknet_leaf_33_clk
rlabel metal2 46536 27440 46536 27440 0 clknet_leaf_34_clk
rlabel metal2 55384 24640 55384 24640 0 clknet_leaf_35_clk
rlabel metal2 48888 12432 48888 12432 0 clknet_leaf_36_clk
rlabel metal2 55272 7560 55272 7560 0 clknet_leaf_37_clk
rlabel metal2 49672 6720 49672 6720 0 clknet_leaf_38_clk
rlabel metal2 45472 12936 45472 12936 0 clknet_leaf_39_clk
rlabel metal2 14952 26264 14952 26264 0 clknet_leaf_3_clk
rlabel metal2 44408 9240 44408 9240 0 clknet_leaf_40_clk
rlabel metal3 30240 7672 30240 7672 0 clknet_leaf_41_clk
rlabel metal2 41720 15960 41720 15960 0 clknet_leaf_42_clk
rlabel metal3 30184 20216 30184 20216 0 clknet_leaf_43_clk
rlabel metal2 27720 22288 27720 22288 0 clknet_leaf_44_clk
rlabel metal2 28168 16968 28168 16968 0 clknet_leaf_45_clk
rlabel metal3 20832 15064 20832 15064 0 clknet_leaf_46_clk
rlabel metal2 29176 12880 29176 12880 0 clknet_leaf_47_clk
rlabel metal2 23240 6384 23240 6384 0 clknet_leaf_48_clk
rlabel metal2 15960 8036 15960 8036 0 clknet_leaf_49_clk
rlabel metal2 14056 19208 14056 19208 0 clknet_leaf_4_clk
rlabel metal3 3080 7560 3080 7560 0 clknet_leaf_50_clk
rlabel metal2 30520 28952 30520 28952 0 clknet_leaf_5_clk
rlabel metal2 21672 31304 21672 31304 0 clknet_leaf_6_clk
rlabel metal2 17248 31864 17248 31864 0 clknet_leaf_7_clk
rlabel metal2 5992 31024 5992 31024 0 clknet_leaf_8_clk
rlabel metal2 5432 36456 5432 36456 0 clknet_leaf_9_clk
rlabel metal3 5600 9016 5600 9016 0 counter10\[0\]
rlabel metal3 12712 16184 12712 16184 0 counter10\[10\]
rlabel metal2 13944 17808 13944 17808 0 counter10\[11\]
rlabel metal2 14224 16296 14224 16296 0 counter10\[12\]
rlabel metal3 13776 15176 13776 15176 0 counter10\[13\]
rlabel metal3 10584 22344 10584 22344 0 counter10\[14\]
rlabel metal2 12712 21672 12712 21672 0 counter10\[15\]
rlabel metal2 11928 21728 11928 21728 0 counter10\[16\]
rlabel metal2 12600 23296 12600 23296 0 counter10\[17\]
rlabel metal2 18536 21784 18536 21784 0 counter10\[18\]
rlabel metal3 17584 19880 17584 19880 0 counter10\[19\]
rlabel metal2 4760 9464 4760 9464 0 counter10\[1\]
rlabel metal2 18088 21224 18088 21224 0 counter10\[20\]
rlabel metal2 16968 19040 16968 19040 0 counter10\[21\]
rlabel metal2 8568 19656 8568 19656 0 counter10\[22\]
rlabel metal2 5544 22792 5544 22792 0 counter10\[23\]
rlabel metal3 5712 19432 5712 19432 0 counter10\[24\]
rlabel metal3 5544 19320 5544 19320 0 counter10\[25\]
rlabel metal3 5040 18424 5040 18424 0 counter10\[26\]
rlabel metal2 8568 17584 8568 17584 0 counter10\[27\]
rlabel metal2 8624 9800 8624 9800 0 counter10\[2\]
rlabel metal2 8680 8372 8680 8372 0 counter10\[3\]
rlabel metal2 11368 7112 11368 7112 0 counter10\[4\]
rlabel metal2 12488 6328 12488 6328 0 counter10\[5\]
rlabel metal2 15288 11312 15288 11312 0 counter10\[6\]
rlabel metal2 13832 12488 13832 12488 0 counter10\[7\]
rlabel metal2 10808 14896 10808 14896 0 counter10\[8\]
rlabel metal3 6608 13608 6608 13608 0 counter10\[9\]
rlabel metal2 44520 47712 44520 47712 0 counter2\[0\]
rlabel metal3 47040 44968 47040 44968 0 counter2\[10\]
rlabel metal2 48104 43988 48104 43988 0 counter2\[11\]
rlabel metal2 49112 43988 49112 43988 0 counter2\[12\]
rlabel metal2 48440 45080 48440 45080 0 counter2\[13\]
rlabel metal2 40712 41496 40712 41496 0 counter2\[14\]
rlabel metal3 42000 42840 42000 42840 0 counter2\[15\]
rlabel metal2 39368 41944 39368 41944 0 counter2\[16\]
rlabel metal2 44520 42224 44520 42224 0 counter2\[17\]
rlabel metal3 41048 45080 41048 45080 0 counter2\[18\]
rlabel metal3 39984 44968 39984 44968 0 counter2\[19\]
rlabel metal2 44072 49784 44072 49784 0 counter2\[1\]
rlabel metal2 43960 45696 43960 45696 0 counter2\[20\]
rlabel metal2 42392 44968 42392 44968 0 counter2\[21\]
rlabel metal2 37128 51240 37128 51240 0 counter2\[22\]
rlabel metal3 37184 47656 37184 47656 0 counter2\[23\]
rlabel metal3 37408 47544 37408 47544 0 counter2\[24\]
rlabel metal2 38248 47824 38248 47824 0 counter2\[25\]
rlabel metal2 43960 49448 43960 49448 0 counter2\[26\]
rlabel metal2 42952 50120 42952 50120 0 counter2\[27\]
rlabel metal3 51800 47544 51800 47544 0 counter2\[2\]
rlabel metal2 52472 48272 52472 48272 0 counter2\[3\]
rlabel metal3 53816 51240 53816 51240 0 counter2\[4\]
rlabel metal2 54040 49392 54040 49392 0 counter2\[5\]
rlabel metal2 53368 44184 53368 44184 0 counter2\[6\]
rlabel metal2 52472 44632 52472 44632 0 counter2\[7\]
rlabel metal2 54152 45416 54152 45416 0 counter2\[8\]
rlabel metal2 55160 44576 55160 44576 0 counter2\[9\]
rlabel metal2 39312 10584 39312 10584 0 counter3\[0\]
rlabel metal2 31080 16800 31080 16800 0 counter3\[10\]
rlabel metal2 33544 18816 33544 18816 0 counter3\[11\]
rlabel metal2 34888 15792 34888 15792 0 counter3\[12\]
rlabel metal2 33992 22568 33992 22568 0 counter3\[13\]
rlabel metal3 34272 23016 34272 23016 0 counter3\[14\]
rlabel metal2 34664 24864 34664 24864 0 counter3\[15\]
rlabel metal2 34440 24752 34440 24752 0 counter3\[16\]
rlabel metal3 30464 27832 30464 27832 0 counter3\[17\]
rlabel metal2 31752 28168 31752 28168 0 counter3\[18\]
rlabel metal2 31416 26880 31416 26880 0 counter3\[19\]
rlabel metal2 39536 10696 39536 10696 0 counter3\[1\]
rlabel metal2 32200 28560 32200 28560 0 counter3\[20\]
rlabel metal3 28280 24024 28280 24024 0 counter3\[21\]
rlabel metal2 28840 22848 28840 22848 0 counter3\[22\]
rlabel metal2 30072 24360 30072 24360 0 counter3\[23\]
rlabel metal2 30520 22064 30520 22064 0 counter3\[24\]
rlabel metal2 31192 20496 31192 20496 0 counter3\[25\]
rlabel metal3 29904 19992 29904 19992 0 counter3\[26\]
rlabel metal2 38304 13608 38304 13608 0 counter3\[27\]
rlabel metal2 40488 6720 40488 6720 0 counter3\[2\]
rlabel metal2 38472 15736 38472 15736 0 counter3\[3\]
rlabel metal3 38304 16184 38304 16184 0 counter3\[4\]
rlabel metal3 37520 20104 37520 20104 0 counter3\[5\]
rlabel metal2 37016 19152 37016 19152 0 counter3\[6\]
rlabel metal3 40432 19320 40432 19320 0 counter3\[7\]
rlabel metal3 38584 19880 38584 19880 0 counter3\[8\]
rlabel metal2 32984 16576 32984 16576 0 counter3\[9\]
rlabel metal2 5992 28560 5992 28560 0 counter4\[0\]
rlabel metal3 25312 26152 25312 26152 0 counter4\[10\]
rlabel metal2 27720 27608 27720 27608 0 counter4\[11\]
rlabel metal2 19208 30352 19208 30352 0 counter4\[12\]
rlabel metal2 20608 32424 20608 32424 0 counter4\[13\]
rlabel metal2 21448 29792 21448 29792 0 counter4\[14\]
rlabel metal2 20440 29344 20440 29344 0 counter4\[15\]
rlabel metal2 20888 23968 20888 23968 0 counter4\[16\]
rlabel metal3 19488 25592 19488 25592 0 counter4\[17\]
rlabel metal3 21280 24584 21280 24584 0 counter4\[18\]
rlabel metal2 20608 25704 20608 25704 0 counter4\[19\]
rlabel metal2 5152 29512 5152 29512 0 counter4\[1\]
rlabel metal2 14728 27328 14728 27328 0 counter4\[20\]
rlabel metal3 13888 27160 13888 27160 0 counter4\[21\]
rlabel metal2 15400 23128 15400 23128 0 counter4\[22\]
rlabel metal3 15456 27272 15456 27272 0 counter4\[23\]
rlabel metal2 16184 31416 16184 31416 0 counter4\[24\]
rlabel metal2 16296 31080 16296 31080 0 counter4\[25\]
rlabel metal2 15960 31444 15960 31444 0 counter4\[26\]
rlabel metal2 15736 31416 15736 31416 0 counter4\[27\]
rlabel metal2 6328 27552 6328 27552 0 counter4\[2\]
rlabel metal2 7336 26320 7336 26320 0 counter4\[3\]
rlabel metal3 25984 32424 25984 32424 0 counter4\[4\]
rlabel metal2 26824 31444 26824 31444 0 counter4\[5\]
rlabel metal2 26768 30744 26768 30744 0 counter4\[6\]
rlabel metal2 26320 30968 26320 30968 0 counter4\[7\]
rlabel metal2 25760 28056 25760 28056 0 counter4\[8\]
rlabel metal3 25424 28840 25424 28840 0 counter4\[9\]
rlabel metal2 54040 39592 54040 39592 0 counter5\[0\]
rlabel metal2 36456 33264 36456 33264 0 counter5\[10\]
rlabel metal3 33656 41384 33656 41384 0 counter5\[11\]
rlabel metal3 34888 41272 34888 41272 0 counter5\[12\]
rlabel metal2 35560 41608 35560 41608 0 counter5\[13\]
rlabel metal2 36568 40712 36568 40712 0 counter5\[14\]
rlabel metal2 31640 37240 31640 37240 0 counter5\[15\]
rlabel metal2 32256 39816 32256 39816 0 counter5\[16\]
rlabel metal2 31528 36288 31528 36288 0 counter5\[17\]
rlabel metal2 32256 33992 32256 33992 0 counter5\[18\]
rlabel metal2 43960 38472 43960 38472 0 counter5\[19\]
rlabel metal3 55384 38136 55384 38136 0 counter5\[1\]
rlabel metal2 44184 39256 44184 39256 0 counter5\[20\]
rlabel metal2 42840 37912 42840 37912 0 counter5\[21\]
rlabel metal2 44632 39536 44632 39536 0 counter5\[22\]
rlabel metal2 42280 36512 42280 36512 0 counter5\[23\]
rlabel metal2 40824 35728 40824 35728 0 counter5\[24\]
rlabel metal2 43400 34944 43400 34944 0 counter5\[25\]
rlabel metal2 41832 35168 41832 35168 0 counter5\[26\]
rlabel metal3 35672 38136 35672 38136 0 counter5\[27\]
rlabel metal3 53144 37352 53144 37352 0 counter5\[2\]
rlabel via2 49000 37240 49000 37240 0 counter5\[3\]
rlabel metal2 49560 39928 49560 39928 0 counter5\[4\]
rlabel metal2 36792 37352 36792 37352 0 counter5\[5\]
rlabel metal3 37128 38136 37128 38136 0 counter5\[6\]
rlabel metal2 35896 33768 35896 33768 0 counter5\[7\]
rlabel metal3 35392 32312 35392 32312 0 counter5\[8\]
rlabel metal2 36568 31388 36568 31388 0 counter5\[9\]
rlabel metal3 27048 7560 27048 7560 0 counter6\[0\]
rlabel metal3 21392 18312 21392 18312 0 counter6\[10\]
rlabel metal2 19376 16184 19376 16184 0 counter6\[11\]
rlabel metal2 22232 17472 22232 17472 0 counter6\[12\]
rlabel metal2 22680 17864 22680 17864 0 counter6\[13\]
rlabel metal2 28112 13160 28112 13160 0 counter6\[14\]
rlabel metal2 27944 13888 27944 13888 0 counter6\[15\]
rlabel metal2 28280 13272 28280 13272 0 counter6\[16\]
rlabel metal3 28784 13160 28784 13160 0 counter6\[17\]
rlabel metal2 32200 10584 32200 10584 0 counter6\[18\]
rlabel metal2 32648 10024 32648 10024 0 counter6\[19\]
rlabel metal2 28000 8344 28000 8344 0 counter6\[1\]
rlabel metal2 32536 11816 32536 11816 0 counter6\[20\]
rlabel metal2 32872 10584 32872 10584 0 counter6\[21\]
rlabel metal2 19544 13888 19544 13888 0 counter6\[22\]
rlabel metal3 18144 13160 18144 13160 0 counter6\[23\]
rlabel metal2 18648 11480 18648 11480 0 counter6\[24\]
rlabel metal2 18760 8372 18760 8372 0 counter6\[25\]
rlabel metal2 22960 12040 22960 12040 0 counter6\[26\]
rlabel metal2 23464 13272 23464 13272 0 counter6\[27\]
rlabel metal2 28168 10584 28168 10584 0 counter6\[2\]
rlabel metal2 26936 8372 26936 8372 0 counter6\[3\]
rlabel metal2 21952 10472 21952 10472 0 counter6\[4\]
rlabel metal2 22120 7392 22120 7392 0 counter6\[5\]
rlabel metal2 24080 19880 24080 19880 0 counter6\[6\]
rlabel metal2 24136 22008 24136 22008 0 counter6\[7\]
rlabel metal3 22624 20888 22624 20888 0 counter6\[8\]
rlabel metal3 24976 20888 24976 20888 0 counter6\[9\]
rlabel metal2 12376 48888 12376 48888 0 counter7\[0\]
rlabel metal2 16632 44044 16632 44044 0 counter7\[10\]
rlabel metal3 14224 42840 14224 42840 0 counter7\[11\]
rlabel metal2 15176 41888 15176 41888 0 counter7\[12\]
rlabel metal3 16800 36568 16800 36568 0 counter7\[13\]
rlabel metal2 16128 35560 16128 35560 0 counter7\[14\]
rlabel metal2 15736 38472 15736 38472 0 counter7\[15\]
rlabel metal2 14728 37576 14728 37576 0 counter7\[16\]
rlabel metal2 7336 35952 7336 35952 0 counter7\[17\]
rlabel metal3 8064 36680 8064 36680 0 counter7\[18\]
rlabel metal3 8568 36568 8568 36568 0 counter7\[19\]
rlabel metal2 12488 49952 12488 49952 0 counter7\[1\]
rlabel metal2 8232 35616 8232 35616 0 counter7\[20\]
rlabel metal2 11312 41272 11312 41272 0 counter7\[21\]
rlabel metal2 10472 39424 10472 39424 0 counter7\[22\]
rlabel metal2 7784 38752 7784 38752 0 counter7\[23\]
rlabel metal2 8904 42896 8904 42896 0 counter7\[24\]
rlabel metal3 9800 43512 9800 43512 0 counter7\[25\]
rlabel metal2 4760 44044 4760 44044 0 counter7\[26\]
rlabel metal2 4816 41272 4816 41272 0 counter7\[27\]
rlabel metal3 13384 48216 13384 48216 0 counter7\[2\]
rlabel metal2 12712 47488 12712 47488 0 counter7\[3\]
rlabel metal2 7896 47040 7896 47040 0 counter7\[4\]
rlabel metal2 7112 49336 7112 49336 0 counter7\[5\]
rlabel metal2 9072 49784 9072 49784 0 counter7\[6\]
rlabel metal3 5208 45976 5208 45976 0 counter7\[7\]
rlabel metal3 5376 41832 5376 41832 0 counter7\[8\]
rlabel metal2 15400 43176 15400 43176 0 counter7\[9\]
rlabel metal3 32032 46536 32032 46536 0 counter8\[0\]
rlabel metal2 23128 38920 23128 38920 0 counter8\[10\]
rlabel metal2 22120 41608 22120 41608 0 counter8\[11\]
rlabel metal2 27496 38360 27496 38360 0 counter8\[12\]
rlabel metal2 27440 36568 27440 36568 0 counter8\[13\]
rlabel metal2 27048 39256 27048 39256 0 counter8\[14\]
rlabel metal3 25984 38808 25984 38808 0 counter8\[15\]
rlabel metal3 21672 35112 21672 35112 0 counter8\[16\]
rlabel metal2 20776 33544 20776 33544 0 counter8\[17\]
rlabel metal2 23016 35336 23016 35336 0 counter8\[18\]
rlabel metal2 22568 34104 22568 34104 0 counter8\[19\]
rlabel metal2 30912 47320 30912 47320 0 counter8\[1\]
rlabel metal2 22344 49448 22344 49448 0 counter8\[20\]
rlabel metal2 22120 49448 22120 49448 0 counter8\[21\]
rlabel metal2 17304 49056 17304 49056 0 counter8\[22\]
rlabel metal3 21336 49112 21336 49112 0 counter8\[23\]
rlabel metal3 21392 45976 21392 45976 0 counter8\[24\]
rlabel metal2 17416 46032 17416 46032 0 counter8\[25\]
rlabel metal3 21672 43400 21672 43400 0 counter8\[26\]
rlabel metal2 22792 45416 22792 45416 0 counter8\[27\]
rlabel metal2 31360 47432 31360 47432 0 counter8\[2\]
rlabel metal2 31080 44688 31080 44688 0 counter8\[3\]
rlabel metal2 26040 45472 26040 45472 0 counter8\[4\]
rlabel metal2 25816 45416 25816 45416 0 counter8\[5\]
rlabel metal2 24696 46312 24696 46312 0 counter8\[6\]
rlabel metal2 24920 49392 24920 49392 0 counter8\[7\]
rlabel metal2 21672 40824 21672 40824 0 counter8\[8\]
rlabel metal3 21280 41272 21280 41272 0 counter8\[9\]
rlabel metal2 47096 23968 47096 23968 0 counter9\[0\]
rlabel metal2 42168 21112 42168 21112 0 counter9\[10\]
rlabel metal3 37856 29288 37856 29288 0 counter9\[11\]
rlabel metal2 38248 28448 38248 28448 0 counter9\[12\]
rlabel metal2 39480 30128 39480 30128 0 counter9\[13\]
rlabel metal2 39704 29848 39704 29848 0 counter9\[14\]
rlabel metal2 40488 24248 40488 24248 0 counter9\[15\]
rlabel metal2 39480 24584 39480 24584 0 counter9\[16\]
rlabel metal3 41440 26152 41440 26152 0 counter9\[17\]
rlabel metal2 42952 25816 42952 25816 0 counter9\[18\]
rlabel metal2 45192 30128 45192 30128 0 counter9\[19\]
rlabel metal3 46200 22232 46200 22232 0 counter9\[1\]
rlabel metal3 44968 29288 44968 29288 0 counter9\[20\]
rlabel metal2 45640 30660 45640 30660 0 counter9\[21\]
rlabel metal2 46312 28112 46312 28112 0 counter9\[22\]
rlabel metal2 49336 31164 49336 31164 0 counter9\[23\]
rlabel metal2 49112 30520 49112 30520 0 counter9\[24\]
rlabel metal3 49056 30296 49056 30296 0 counter9\[25\]
rlabel metal2 52472 30632 52472 30632 0 counter9\[26\]
rlabel metal2 41384 22288 41384 22288 0 counter9\[27\]
rlabel metal2 45640 22736 45640 22736 0 counter9\[2\]
rlabel metal2 45976 21560 45976 21560 0 counter9\[3\]
rlabel metal2 50456 22008 50456 22008 0 counter9\[4\]
rlabel metal3 52304 23128 52304 23128 0 counter9\[5\]
rlabel metal2 51184 24696 51184 24696 0 counter9\[6\]
rlabel metal2 52584 27160 52584 27160 0 counter9\[7\]
rlabel metal2 49280 27160 49280 27160 0 counter9\[8\]
rlabel metal2 40824 22512 40824 22512 0 counter9\[9\]
rlabel metal3 52192 11592 52192 11592 0 counter\[0\]
rlabel metal3 45080 15288 45080 15288 0 counter\[10\]
rlabel metal2 46032 15288 46032 15288 0 counter\[11\]
rlabel metal2 46312 16520 46312 16520 0 counter\[12\]
rlabel metal2 53368 14392 53368 14392 0 counter\[13\]
rlabel metal2 53144 14168 53144 14168 0 counter\[14\]
rlabel metal3 53200 13720 53200 13720 0 counter\[15\]
rlabel metal2 53816 14168 53816 14168 0 counter\[16\]
rlabel metal3 52528 18200 52528 18200 0 counter\[17\]
rlabel metal2 52472 18368 52472 18368 0 counter\[18\]
rlabel metal2 53536 18424 53536 18424 0 counter\[19\]
rlabel metal3 52360 11480 52360 11480 0 counter\[1\]
rlabel metal2 53816 17976 53816 17976 0 counter\[20\]
rlabel metal2 51912 8288 51912 8288 0 counter\[21\]
rlabel metal2 49112 6720 49112 6720 0 counter\[22\]
rlabel metal2 52584 6832 52584 6832 0 counter\[23\]
rlabel metal3 52976 7336 52976 7336 0 counter\[24\]
rlabel metal2 52472 10024 52472 10024 0 counter\[25\]
rlabel metal2 53480 10640 53480 10640 0 counter\[26\]
rlabel metal3 45136 11592 45136 11592 0 counter\[27\]
rlabel metal2 45864 12320 45864 12320 0 counter\[2\]
rlabel metal2 46088 11704 46088 11704 0 counter\[3\]
rlabel metal2 45976 11368 45976 11368 0 counter\[4\]
rlabel metal2 43960 10248 43960 10248 0 counter\[5\]
rlabel metal2 44744 9632 44744 9632 0 counter\[6\]
rlabel metal2 45528 10136 45528 10136 0 counter\[7\]
rlabel metal2 45640 9912 45640 9912 0 counter\[8\]
rlabel metal2 45864 15736 45864 15736 0 counter\[9\]
rlabel metal2 55384 5320 55384 5320 0 cout1
rlabel metal2 56 2198 56 2198 0 cout10
rlabel metal2 50008 56280 50008 56280 0 cout2
rlabel metal2 43736 2198 43736 2198 0 cout3
rlabel metal3 1638 21560 1638 21560 0 cout4
rlabel metal2 55384 49392 55384 49392 0 cout5
rlabel metal2 21560 2198 21560 2198 0 cout6
rlabel metal2 6440 56280 6440 56280 0 cout7
rlabel metal2 27832 56280 27832 56280 0 cout8
rlabel metal3 57330 26936 57330 26936 0 cout9
rlabel metal2 56280 5432 56280 5432 0 net1
rlabel metal2 56448 26264 56448 26264 0 net10
rlabel metal2 34832 50456 34832 50456 0 net100
rlabel metal2 39144 47712 39144 47712 0 net101
rlabel metal3 41328 45304 41328 45304 0 net102
rlabel metal2 36232 44576 36232 44576 0 net103
rlabel metal2 38360 46368 38360 46368 0 net104
rlabel metal2 42392 43876 42392 43876 0 net105
rlabel metal2 37240 42280 37240 42280 0 net106
rlabel metal2 39480 43232 39480 43232 0 net107
rlabel metal2 38584 40712 38584 40712 0 net108
rlabel metal2 46368 44184 46368 44184 0 net109
rlabel metal2 20720 45192 20720 45192 0 net11
rlabel metal3 49784 43736 49784 43736 0 net110
rlabel metal2 45864 43876 45864 43876 0 net111
rlabel metal2 44576 44184 44576 44184 0 net112
rlabel metal2 53816 45416 53816 45416 0 net113
rlabel metal2 52080 45752 52080 45752 0 net114
rlabel metal2 50344 45416 50344 45416 0 net115
rlabel metal2 50792 42056 50792 42056 0 net116
rlabel metal2 52080 47320 52080 47320 0 net117
rlabel metal2 50344 50848 50344 50848 0 net118
rlabel metal3 49672 48888 49672 48888 0 net119
rlabel metal2 19320 43876 19320 43876 0 net12
rlabel metal2 48048 47544 48048 47544 0 net120
rlabel metal2 36288 13832 36288 13832 0 net121
rlabel metal2 26712 20440 26712 20440 0 net122
rlabel metal2 29848 20440 29848 20440 0 net123
rlabel metal2 28448 21672 28448 21672 0 net124
rlabel metal2 28224 24808 28224 24808 0 net125
rlabel metal2 26712 23072 26712 23072 0 net126
rlabel metal3 25200 24024 25200 24024 0 net127
rlabel metal2 30744 29736 30744 29736 0 net128
rlabel metal2 29288 27384 29288 27384 0 net129
rlabel metal3 16520 45304 16520 45304 0 net13
rlabel metal2 30072 30464 30072 30464 0 net130
rlabel metal2 27272 29736 27272 29736 0 net131
rlabel metal2 33768 26712 33768 26712 0 net132
rlabel metal2 32200 25984 32200 25984 0 net133
rlabel metal3 35224 22232 35224 22232 0 net134
rlabel metal2 31864 23072 31864 23072 0 net135
rlabel metal2 32760 15232 32760 15232 0 net136
rlabel metal2 31640 18872 31640 18872 0 net137
rlabel metal2 29064 16856 29064 16856 0 net138
rlabel metal2 30856 16296 30856 16296 0 net139
rlabel metal2 18760 46592 18760 46592 0 net14
rlabel metal3 36624 20552 36624 20552 0 net140
rlabel metal2 38864 18648 38864 18648 0 net141
rlabel metal2 35112 17920 35112 17920 0 net142
rlabel metal2 34384 20216 34384 20216 0 net143
rlabel metal3 40376 16184 40376 16184 0 net144
rlabel metal2 36400 15400 36400 15400 0 net145
rlabel metal2 16520 33824 16520 33824 0 net146
rlabel metal2 13664 32648 13664 32648 0 net147
rlabel metal2 10808 31892 10808 31892 0 net148
rlabel metal2 13944 30856 13944 30856 0 net149
rlabel metal2 18704 48440 18704 48440 0 net15
rlabel metal2 13776 27944 13776 27944 0 net150
rlabel metal3 13608 23240 13608 23240 0 net151
rlabel metal2 11480 26824 11480 26824 0 net152
rlabel metal2 10808 29120 10808 29120 0 net153
rlabel metal2 18536 26600 18536 26600 0 net154
rlabel metal2 19600 24808 19600 24808 0 net155
rlabel metal3 17136 24920 17136 24920 0 net156
rlabel metal2 18872 22456 18872 22456 0 net157
rlabel metal2 17416 29120 17416 29120 0 net158
rlabel metal2 19320 30520 19320 30520 0 net159
rlabel metal2 15176 49504 15176 49504 0 net16
rlabel metal2 18312 31780 18312 31780 0 net160
rlabel metal2 17752 29848 17752 29848 0 net161
rlabel metal2 25592 27776 25592 27776 0 net162
rlabel metal2 22456 27944 22456 27944 0 net163
rlabel metal2 22792 29736 22792 29736 0 net164
rlabel metal2 23016 26208 23016 26208 0 net165
rlabel metal2 28392 32872 28392 32872 0 net166
rlabel metal2 24808 30856 24808 30856 0 net167
rlabel metal2 24472 34048 24472 34048 0 net168
rlabel metal2 22792 32872 22792 32872 0 net169
rlabel metal2 19320 51688 19320 51688 0 net17
rlabel metal3 33264 38920 33264 38920 0 net170
rlabel metal2 43960 35616 43960 35616 0 net171
rlabel metal2 41272 33824 41272 33824 0 net172
rlabel metal2 38920 34552 38920 34552 0 net173
rlabel metal2 40376 36120 40376 36120 0 net174
rlabel metal2 45640 39872 45640 39872 0 net175
rlabel metal2 44968 37576 44968 37576 0 net176
rlabel metal2 41944 39256 41944 39256 0 net177
rlabel metal2 41832 38528 41832 38528 0 net178
rlabel metal2 30128 34216 30128 34216 0 net179
rlabel metal2 20776 50120 20776 50120 0 net18
rlabel metal2 29400 36008 29400 36008 0 net180
rlabel metal2 30408 38696 30408 38696 0 net181
rlabel metal2 29624 38276 29624 38276 0 net182
rlabel metal2 34384 40488 34384 40488 0 net183
rlabel metal2 34440 43456 34440 43456 0 net184
rlabel metal2 32312 41664 32312 41664 0 net185
rlabel metal2 30184 41440 30184 41440 0 net186
rlabel metal3 37016 34216 37016 34216 0 net187
rlabel metal2 34104 30464 34104 30464 0 net188
rlabel metal2 32704 31752 32704 31752 0 net189
rlabel metal2 21672 33600 21672 33600 0 net19
rlabel metal2 33824 34328 33824 34328 0 net190
rlabel metal2 39704 38360 39704 38360 0 net191
rlabel metal3 35112 37352 35112 37352 0 net192
rlabel metal2 21336 14056 21336 14056 0 net193
rlabel metal2 20776 12488 20776 12488 0 net194
rlabel metal2 16688 8344 16688 8344 0 net195
rlabel metal2 16520 11312 16520 11312 0 net196
rlabel metal3 15232 12824 15232 12824 0 net197
rlabel metal2 17864 14168 17864 14168 0 net198
rlabel metal3 34776 12376 34776 12376 0 net199
rlabel metal2 1848 4648 1848 4648 0 net2
rlabel metal2 21952 35784 21952 35784 0 net20
rlabel metal2 30744 13664 30744 13664 0 net200
rlabel metal2 30744 9464 30744 9464 0 net201
rlabel metal2 30016 12264 30016 12264 0 net202
rlabel metal2 26936 15624 26936 15624 0 net203
rlabel metal2 26488 17920 26488 17920 0 net204
rlabel metal3 23184 15848 23184 15848 0 net205
rlabel metal2 26040 14168 26040 14168 0 net206
rlabel metal2 24808 18144 24808 18144 0 net207
rlabel metal2 20160 16968 20160 16968 0 net208
rlabel metal2 17304 16576 17304 16576 0 net209
rlabel metal2 18648 34608 18648 34608 0 net21
rlabel metal2 18872 17920 18872 17920 0 net210
rlabel metal2 23240 21280 23240 21280 0 net211
rlabel metal3 19152 20216 19152 20216 0 net212
rlabel metal2 22400 21784 22400 21784 0 net213
rlabel metal2 21952 20104 21952 20104 0 net214
rlabel metal2 2688 41272 2688 41272 0 net215
rlabel metal2 2688 44408 2688 44408 0 net216
rlabel metal2 7280 44408 7280 44408 0 net217
rlabel metal2 6832 42168 6832 42168 0 net218
rlabel metal2 5656 39704 5656 39704 0 net219
rlabel metal2 19712 35896 19712 35896 0 net22
rlabel metal2 8568 39256 8568 39256 0 net220
rlabel metal2 9800 40824 9800 40824 0 net221
rlabel metal2 7112 33600 7112 33600 0 net222
rlabel metal2 11256 36736 11256 36736 0 net223
rlabel metal2 6440 36736 6440 36736 0 net224
rlabel metal2 5208 35504 5208 35504 0 net225
rlabel metal2 12600 38136 12600 38136 0 net226
rlabel metal2 13608 39144 13608 39144 0 net227
rlabel metal2 14000 35784 14000 35784 0 net228
rlabel metal2 15288 36960 15288 36960 0 net229
rlabel metal2 23016 40096 23016 40096 0 net23
rlabel metal3 13384 40488 13384 40488 0 net230
rlabel metal3 11312 41048 11312 41048 0 net231
rlabel metal2 13888 43736 13888 43736 0 net232
rlabel metal3 17024 42168 17024 42168 0 net233
rlabel metal2 2856 43232 2856 43232 0 net234
rlabel metal3 3192 45976 3192 45976 0 net235
rlabel metal2 27832 39928 27832 39928 0 net24
rlabel metal3 25144 36568 25144 36568 0 net25
rlabel metal2 25368 38528 25368 38528 0 net26
rlabel metal2 20216 42280 20216 42280 0 net27
rlabel metal2 20944 38920 20944 38920 0 net28
rlabel metal2 18088 40824 18088 40824 0 net29
rlabel metal2 48776 53340 48776 53340 0 net3
rlabel metal2 17920 39032 17920 39032 0 net30
rlabel metal2 38696 23464 38696 23464 0 net31
rlabel metal2 50344 31500 50344 31500 0 net32
rlabel metal2 46480 29624 46480 29624 0 net33
rlabel metal2 46648 31500 46648 31500 0 net34
rlabel metal3 47320 34328 47320 34328 0 net35
rlabel metal2 44240 27944 44240 27944 0 net36
rlabel metal2 43848 31752 43848 31752 0 net37
rlabel metal2 42336 28504 42336 28504 0 net38
rlabel metal2 43512 30464 43512 30464 0 net39
rlabel metal2 43400 4368 43400 4368 0 net4
rlabel metal2 40880 25592 40880 25592 0 net40
rlabel metal2 38696 27776 38696 27776 0 net41
rlabel metal2 37016 24864 37016 24864 0 net42
rlabel metal2 38360 24752 38360 24752 0 net43
rlabel metal2 38360 31892 38360 31892 0 net44
rlabel metal3 37352 31080 37352 31080 0 net45
rlabel metal2 36120 28168 36120 28168 0 net46
rlabel metal2 34440 28672 34440 28672 0 net47
rlabel metal3 40320 20216 40320 20216 0 net48
rlabel metal2 38752 22456 38752 22456 0 net49
rlabel metal2 1848 22008 1848 22008 0 net5
rlabel metal2 6496 16968 6496 16968 0 net50
rlabel metal2 4424 15960 4424 15960 0 net51
rlabel metal3 3360 20552 3360 20552 0 net52
rlabel metal2 3192 20356 3192 20356 0 net53
rlabel metal2 3472 23240 3472 23240 0 net54
rlabel metal2 6496 20104 6496 20104 0 net55
rlabel metal2 15512 19432 15512 19432 0 net56
rlabel metal3 15680 22456 15680 22456 0 net57
rlabel metal2 14784 20104 14784 20104 0 net58
rlabel metal3 13720 23800 13720 23800 0 net59
rlabel metal2 56504 49448 56504 49448 0 net6
rlabel metal2 10360 23576 10360 23576 0 net60
rlabel metal2 9856 20216 9856 20216 0 net61
rlabel metal2 10640 20216 10640 20216 0 net62
rlabel metal2 7336 22400 7336 22400 0 net63
rlabel metal2 15064 16184 15064 16184 0 net64
rlabel metal2 12208 15960 12208 15960 0 net65
rlabel metal2 10696 18872 10696 18872 0 net66
rlabel metal2 9632 16184 9632 16184 0 net67
rlabel metal2 42336 12264 42336 12264 0 net68
rlabel metal2 54936 10528 54936 10528 0 net69
rlabel metal2 22008 4648 22008 4648 0 net7
rlabel metal2 50344 9632 50344 9632 0 net70
rlabel metal3 54936 7560 54936 7560 0 net71
rlabel metal2 50456 7168 50456 7168 0 net72
rlabel metal2 46984 7336 46984 7336 0 net73
rlabel metal3 49280 8232 49280 8232 0 net74
rlabel metal2 54824 18144 54824 18144 0 net75
rlabel metal3 54152 19096 54152 19096 0 net76
rlabel metal2 50344 19264 50344 19264 0 net77
rlabel metal3 50120 20216 50120 20216 0 net78
rlabel metal2 54152 15008 54152 15008 0 net79
rlabel metal3 3584 50680 3584 50680 0 net8
rlabel metal3 52024 15960 52024 15960 0 net80
rlabel metal2 48216 15008 48216 15008 0 net81
rlabel metal3 49784 15400 49784 15400 0 net82
rlabel metal3 47096 17752 47096 17752 0 net83
rlabel metal2 43736 19264 43736 19264 0 net84
rlabel metal3 41720 17528 41720 17528 0 net85
rlabel metal3 45864 15960 45864 15960 0 net86
rlabel metal3 47152 9912 47152 9912 0 net87
rlabel metal2 45528 7784 45528 7784 0 net88
rlabel metal2 42616 9912 42616 9912 0 net89
rlabel metal2 27272 53368 27272 53368 0 net9
rlabel metal2 41832 10304 41832 10304 0 net90
rlabel metal2 47656 12656 47656 12656 0 net91
rlabel metal3 45192 12824 45192 12824 0 net92
rlabel metal2 39816 13440 39816 13440 0 net93
rlabel metal2 48944 11480 48944 11480 0 net94
rlabel metal2 40824 51072 40824 51072 0 net95
rlabel metal2 41776 49112 41776 49112 0 net96
rlabel metal2 39704 49728 39704 49728 0 net97
rlabel metal2 34664 48160 34664 48160 0 net98
rlabel metal2 34440 48552 34440 48552 0 net99
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
